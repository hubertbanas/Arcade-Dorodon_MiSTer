library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_cpu1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_cpu1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"B3",X"00",X"25",X"9F",X"DE",X"00",X"B0",X"DE",X"00",X"C0",X"25",X"BF",X"DE",
		X"00",X"B0",X"DE",X"00",X"C0",X"25",X"DF",X"DE",X"00",X"B0",X"DE",X"00",X"C0",X"25",X"FF",X"DE",
		X"00",X"B0",X"DE",X"00",X"C0",X"89",X"DE",X"76",X"00",X"62",X"B3",X"00",X"71",X"00",X"C0",X"89",
		X"FB",X"7A",X"00",X"01",X"FF",X"FF",X"FF",X"FF",X"7A",X"9E",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7A",X"34",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"4B",X"27",X"60",X"5C",X"7A",X"9B",X"3B",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"59",X"FF",X"67",X"B6",X"0D",X"E3",X"4B",X"00",X"80",X"A4",X"6E",X"17",X"A4",X"D4",X"1A",X"A4",
		X"06",X"2B",X"A4",X"BA",X"1A",X"A4",X"55",X"17",X"A4",X"C6",X"02",X"59",X"FF",X"67",X"EE",X"DE",
		X"00",X"A0",X"A4",X"BA",X"1A",X"A4",X"A2",X"5B",X"1A",X"1C",X"00",X"B3",X"03",X"CB",X"EE",X"A4",
		X"71",X"4C",X"B3",X"20",X"A4",X"A9",X"4D",X"25",X"01",X"A4",X"71",X"4C",X"B3",X"20",X"A4",X"A9",
		X"4D",X"DC",X"89",X"E9",X"B5",X"00",X"A4",X"60",X"4C",X"A4",X"2B",X"01",X"76",X"02",X"90",X"19",
		X"86",X"9B",X"8C",X"01",X"A4",X"99",X"4C",X"76",X"5F",X"60",X"19",X"6D",X"76",X"F8",X"0E",X"37",
		X"D8",X"61",X"A4",X"36",X"1F",X"DE",X"66",X"60",X"EE",X"DE",X"67",X"60",X"DE",X"65",X"60",X"DE",
		X"6E",X"60",X"DE",X"6F",X"60",X"7A",X"F7",X"03",X"76",X"1C",X"60",X"EE",X"F8",X"76",X"21",X"60",
		X"F8",X"A4",X"CD",X"3C",X"76",X"5F",X"60",X"19",X"CD",X"7A",X"1B",X"01",X"25",X"09",X"DE",X"5E",
		X"60",X"7A",X"5F",X"03",X"CB",X"97",X"B3",X"1F",X"A4",X"28",X"05",X"01",X"DC",X"B5",X"97",X"66",
		X"CB",X"4B",X"CD",X"61",X"F4",X"00",X"F3",X"2B",X"02",X"4B",X"5B",X"60",X"F4",X"00",X"F3",X"2B",
		X"02",X"25",X"03",X"DE",X"5B",X"60",X"25",X"FF",X"76",X"03",X"90",X"B6",X"E9",X"8B",X"76",X"E2",
		X"0B",X"19",X"99",X"04",X"B3",X"00",X"D6",X"26",X"51",X"19",X"8E",X"76",X"30",X"68",X"D6",X"D1",
		X"7B",X"21",X"9B",X"D9",X"01",X"D3",X"7A",X"26",X"02",X"71",X"00",X"C7",X"7B",X"D3",X"7A",X"FC",
		X"01",X"4B",X"0C",X"62",X"19",X"04",X"9B",X"8B",X"08",X"19",X"75",X"DE",X"0C",X"62",X"19",X"4A",
		X"76",X"FF",X"FF",X"F2",X"01",X"A4",X"2C",X"3C",X"7A",X"77",X"02",X"00",X"76",X"5E",X"60",X"03",
		X"F8",X"72",X"4B",X"21",X"D3",X"F4",X"1D",X"ED",X"08",X"65",X"F4",X"0A",X"EA",X"03",X"DE",X"61",
		X"D3",X"4B",X"5F",X"60",X"19",X"72",X"ED",X"0E",X"76",X"08",X"00",X"8E",X"A9",X"F7",X"5F",X"03",
		X"CB",X"76",X"FA",X"FF",X"8E",X"A9",X"76",X"01",X"60",X"19",X"6D",X"4B",X"00",X"80",X"0E",X"DC",
		X"3E",X"01",X"B6",X"47",X"97",X"66",X"CB",X"4B",X"CD",X"61",X"F4",X"00",X"F3",X"C1",X"02",X"4B",
		X"5B",X"60",X"F4",X"00",X"F3",X"C1",X"02",X"25",X"03",X"DE",X"5B",X"60",X"25",X"FF",X"76",X"03",
		X"90",X"B6",X"EB",X"8B",X"76",X"E2",X"0B",X"19",X"99",X"04",X"B3",X"00",X"D6",X"26",X"51",X"19",
		X"8E",X"76",X"30",X"68",X"D6",X"D1",X"7B",X"21",X"9B",X"6F",X"02",X"D3",X"7A",X"BC",X"02",X"71",
		X"00",X"C7",X"7B",X"D3",X"7A",X"92",X"02",X"A4",X"BD",X"3D",X"66",X"76",X"01",X"60",X"19",X"F4",
		X"3E",X"7A",X"84",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"76",X"5E",X"60",X"03",X"F8",X"72",X"4B",X"21",X"D3",X"F4",X"1D",X"ED",X"08",X"65",
		X"F4",X"0A",X"EA",X"03",X"DE",X"61",X"D3",X"4B",X"5F",X"60",X"19",X"72",X"ED",X"0E",X"76",X"08",
		X"00",X"8E",X"A9",X"F7",X"5F",X"03",X"CB",X"76",X"FA",X"FF",X"8E",X"A9",X"76",X"01",X"60",X"19",
		X"6D",X"DC",X"3E",X"01",X"B6",X"43",X"EE",X"DE",X"5B",X"60",X"DE",X"00",X"A0",X"DE",X"C9",X"61",
		X"A4",X"24",X"50",X"DE",X"CD",X"61",X"DE",X"5E",X"60",X"7A",X"57",X"49",X"A4",X"F9",X"02",X"A4",
		X"12",X"03",X"EE",X"76",X"68",X"60",X"F8",X"C0",X"F8",X"C0",X"F8",X"76",X"00",X"60",X"B3",X"1C",
		X"F8",X"C0",X"89",X"FC",X"A4",X"2F",X"03",X"0E",X"B5",X"B3",X"09",X"76",X"73",X"60",X"EE",X"5C",
		X"F8",X"EE",X"C0",X"F8",X"C0",X"F8",X"C0",X"89",X"F6",X"B5",X"A4",X"FB",X"5B",X"A4",X"BA",X"1A",
		X"B5",X"00",X"76",X"80",X"D3",X"B3",X"09",X"CB",X"D9",X"76",X"02",X"2F",X"B3",X"07",X"D9",X"22",
		X"00",X"D9",X"C0",X"F8",X"C0",X"89",X"F7",X"25",X"FF",X"F8",X"C0",X"DC",X"89",X"E9",X"B5",X"B3",
		X"32",X"EE",X"76",X"1C",X"60",X"F8",X"C0",X"89",X"FC",X"B5",X"97",X"4B",X"5B",X"60",X"F4",X"00",
		X"7D",X"04",X"5E",X"DE",X"5B",X"60",X"4B",X"CD",X"61",X"F4",X"00",X"7D",X"01",X"5E",X"DE",X"CD",
		X"61",X"4B",X"00",X"90",X"19",X"B8",X"ED",X"05",X"25",X"05",X"DE",X"CD",X"61",X"01",X"B5",X"76",
		X"5F",X"60",X"19",X"5A",X"19",X"CD",X"76",X"1C",X"60",X"EE",X"F8",X"76",X"21",X"60",X"F8",X"A4",
		X"CD",X"3C",X"EE",X"DE",X"00",X"A0",X"A4",X"25",X"25",X"25",X"01",X"DE",X"E2",X"61",X"EE",X"DE",
		X"C8",X"61",X"F7",X"01",X"00",X"76",X"00",X"90",X"19",X"24",X"7D",X"27",X"4B",X"5E",X"60",X"F4",
		X"02",X"2C",X"04",X"19",X"86",X"7D",X"34",X"CB",X"A4",X"A5",X"1C",X"A4",X"E5",X"27",X"A4",X"55",
		X"27",X"A4",X"5A",X"2D",X"B3",X"01",X"A4",X"2D",X"01",X"DC",X"89",X"D9",X"1A",X"D4",X"00",X"00",
		X"00",X"00",X"00",X"4B",X"5F",X"60",X"19",X"10",X"DE",X"5F",X"60",X"A4",X"36",X"1F",X"DE",X"66",
		X"60",X"EE",X"DE",X"67",X"60",X"76",X"5E",X"60",X"9E",X"1A",X"16",X"4B",X"5F",X"60",X"19",X"9C",
		X"DE",X"5F",X"60",X"A4",X"36",X"1F",X"DE",X"66",X"60",X"DE",X"67",X"60",X"7A",X"60",X"49",X"9E",
		X"9E",X"EE",X"7A",X"6C",X"49",X"76",X"68",X"60",X"F8",X"C0",X"F8",X"C0",X"F8",X"C0",X"F8",X"C0",
		X"F8",X"C0",X"F8",X"C0",X"F8",X"C0",X"F8",X"25",X"FF",X"76",X"9D",X"60",X"B3",X"06",X"F8",X"C0",
		X"89",X"FC",X"EE",X"DE",X"9F",X"60",X"DE",X"A2",X"60",X"76",X"1C",X"D6",X"37",X"63",X"60",X"76",
		X"5F",X"60",X"19",X"AC",X"A4",X"0A",X"03",X"A4",X"E5",X"1B",X"EE",X"DE",X"60",X"60",X"8B",X"DE",
		X"62",X"60",X"25",X"0C",X"DE",X"61",X"60",X"A4",X"C6",X"1C",X"A4",X"44",X"21",X"A4",X"BC",X"5D",
		X"A4",X"64",X"1D",X"A4",X"77",X"1D",X"A4",X"D1",X"1D",X"A4",X"8B",X"1E",X"B3",X"08",X"25",X"05",
		X"76",X"E1",X"D4",X"A4",X"7D",X"1E",X"A4",X"E0",X"1E",X"A4",X"26",X"28",X"B3",X"05",X"25",X"05",
		X"76",X"E1",X"D4",X"A4",X"7D",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D9",
		X"76",X"1C",X"60",X"D9",X"71",X"00",X"82",X"D9",X"71",X"01",X"06",X"D9",X"71",X"02",X"0F",X"A4",
		X"7F",X"1F",X"D9",X"F8",X"03",X"D9",X"A3",X"04",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"D9",X"71",
		X"00",X"81",X"7A",X"D5",X"04",X"D9",X"76",X"70",X"60",X"B6",X"57",X"D4",X"00",X"3D",X"19",X"15",
		X"D9",X"08",X"00",X"B6",X"57",X"6D",X"07",X"3D",X"54",X"02",X"F4",X"05",X"ED",X"0A",X"4B",X"E2",
		X"61",X"F4",X"00",X"25",X"05",X"ED",X"01",X"5C",X"D9",X"F8",X"01",X"B6",X"57",X"3D",X"6D",X"03",
		X"3D",X"54",X"07",X"F4",X"08",X"ED",X"1A",X"72",X"A4",X"36",X"1F",X"5C",X"04",X"4B",X"65",X"60",
		X"F4",X"00",X"7D",X"05",X"4B",X"67",X"60",X"1A",X"03",X"4B",X"66",X"60",X"67",X"65",X"2C",X"01",
		X"5C",X"D9",X"F8",X"02",X"B5",X"EE",X"DE",X"C9",X"61",X"A4",X"CF",X"33",X"A4",X"77",X"1D",X"A4",
		X"85",X"04",X"A4",X"FE",X"28",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"25",X"81",X"DE",X"21",X"60",
		X"A4",X"F4",X"30",X"A4",X"1C",X"31",X"A4",X"54",X"31",X"A4",X"77",X"1D",X"A4",X"F4",X"1E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"76",X"1F",X"60",X"A4",X"7F",X"1F",X"F8",X"C0",X"A3",X"A4",X"C7",
		X"1F",X"A4",X"8F",X"17",X"B3",X"B4",X"A4",X"28",X"05",X"A4",X"C1",X"2A",X"EE",X"DE",X"21",X"60",
		X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"1A",X"19",X"76",X"01",X"90",X"A4",X"5A",X"2D",X"19",X"22",
		X"7D",X"FC",X"19",X"22",X"ED",X"FC",X"CB",X"A4",X"3A",X"03",X"A4",X"8F",X"17",X"DC",X"89",X"E8",
		X"B5",X"A4",X"44",X"21",X"A4",X"E3",X"33",X"00",X"00",X"00",X"A4",X"92",X"31",X"A4",X"DA",X"30",
		X"A4",X"CF",X"30",X"A4",X"44",X"31",X"25",X"03",X"DE",X"9B",X"61",X"A4",X"15",X"2B",X"A4",X"F4",
		X"30",X"A4",X"1C",X"31",X"A4",X"54",X"31",X"A4",X"F4",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",
		X"D9",X"76",X"1C",X"60",X"D9",X"71",X"00",X"82",X"D9",X"71",X"01",X"06",X"D9",X"71",X"02",X"0F",
		X"A4",X"7F",X"1F",X"D9",X"F8",X"03",X"D9",X"A3",X"04",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"D9",
		X"71",X"00",X"81",X"76",X"1C",X"D6",X"37",X"63",X"60",X"EE",X"DE",X"60",X"60",X"8B",X"DE",X"62",
		X"60",X"25",X"0C",X"DE",X"61",X"60",X"A4",X"C6",X"1C",X"A4",X"AE",X"05",X"1A",X"23",X"15",X"05",
		X"00",X"76",X"2B",X"60",X"D4",X"00",X"22",X"6D",X"03",X"7D",X"08",X"40",X"77",X"F4",X"04",X"ED",
		X"F5",X"1A",X"0D",X"A4",X"61",X"30",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"D9",X"71",X"00",X"81",
		X"B5",X"4B",X"65",X"60",X"F4",X"00",X"7D",X"05",X"76",X"67",X"60",X"1A",X"03",X"76",X"66",X"60",
		X"9E",X"22",X"97",X"A4",X"77",X"1D",X"01",X"D9",X"76",X"26",X"60",X"D9",X"71",X"00",X"82",X"D9",
		X"71",X"01",X"58",X"D9",X"71",X"02",X"56",X"EE",X"D9",X"F8",X"03",X"D9",X"F8",X"04",X"76",X"00",
		X"60",X"19",X"FE",X"25",X"FF",X"A4",X"4C",X"1E",X"7A",X"30",X"07",X"A4",X"C1",X"2A",X"EE",X"DE",
		X"C9",X"61",X"A4",X"4C",X"1E",X"7A",X"41",X"05",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"A4",X"CF",X"33",X"76",X"66",X"60",X"4B",X"65",X"60",X"F4",X"00",X"7D",X"03",X"76",
		X"67",X"60",X"D1",X"D1",X"66",X"A4",X"85",X"04",X"3E",X"9E",X"9E",X"A4",X"FE",X"28",X"A4",X"C7",
		X"1F",X"A4",X"8F",X"17",X"25",X"81",X"DE",X"21",X"60",X"A4",X"F4",X"30",X"A4",X"1C",X"31",X"A4",
		X"54",X"31",X"A4",X"77",X"1D",X"A4",X"F4",X"1E",X"76",X"01",X"D1",X"00",X"00",X"00",X"76",X"1F",
		X"60",X"A4",X"7F",X"1F",X"F8",X"C0",X"A3",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"B3",X"B4",X"A4",
		X"28",X"05",X"A4",X"1B",X"0A",X"EE",X"DE",X"21",X"60",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"A4",
		X"44",X"21",X"A4",X"E3",X"33",X"00",X"00",X"00",X"A4",X"92",X"31",X"A4",X"44",X"31",X"A4",X"54",
		X"31",X"A4",X"DA",X"30",X"A4",X"CF",X"30",X"A4",X"15",X"2B",X"EE",X"DE",X"60",X"60",X"8B",X"DE",
		X"62",X"60",X"25",X"0C",X"DE",X"61",X"60",X"A4",X"C6",X"1C",X"76",X"1C",X"D6",X"37",X"63",X"60",
		X"A4",X"F4",X"1E",X"76",X"01",X"D1",X"00",X"00",X"00",X"D9",X"76",X"1C",X"60",X"D9",X"71",X"00",
		X"82",X"D9",X"71",X"01",X"06",X"D9",X"71",X"02",X"0F",X"A4",X"7F",X"1F",X"D9",X"F8",X"03",X"D9",
		X"A3",X"04",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"D9",X"71",X"00",X"81",X"A4",X"AE",X"05",X"76",
		X"26",X"60",X"71",X"82",X"C0",X"71",X"58",X"C0",X"71",X"56",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",
		X"A4",X"E3",X"35",X"D9",X"76",X"B6",X"61",X"D9",X"71",X"00",X"60",X"D9",X"71",X"01",X"00",X"D9",
		X"71",X"02",X"00",X"D9",X"71",X"03",X"B4",X"EE",X"DE",X"B5",X"61",X"DE",X"B4",X"61",X"DE",X"E1",
		X"61",X"76",X"CE",X"61",X"B3",X"05",X"EE",X"F8",X"C0",X"89",X"FC",X"76",X"5F",X"60",X"19",X"F4",
		X"76",X"96",X"61",X"71",X"58",X"C0",X"71",X"56",X"C0",X"71",X"08",X"25",X"08",X"DE",X"98",X"61",
		X"15",X"00",X"00",X"B6",X"2F",X"99",X"61",X"76",X"5F",X"60",X"19",X"11",X"A4",X"FD",X"45",X"A4",
		X"3A",X"46",X"1A",X"06",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"A4",X"5A",X"2D",X"76",X"5F",X"60",
		X"19",X"05",X"ED",X"08",X"76",X"02",X"90",X"19",X"69",X"9B",X"5E",X"09",X"A4",X"B1",X"39",X"A4",
		X"6D",X"2B",X"4B",X"E1",X"61",X"F4",X"00",X"ED",X"03",X"A4",X"7E",X"40",X"A4",X"37",X"5F",X"A4",
		X"FF",X"35",X"A4",X"99",X"3A",X"B3",X"04",X"7A",X"60",X"21",X"15",X"05",X"00",X"19",X"FA",X"F3",
		X"C8",X"07",X"40",X"89",X"F8",X"7A",X"EE",X"07",X"66",X"C0",X"C0",X"4B",X"28",X"60",X"AC",X"EA",
		X"02",X"B6",X"CF",X"F4",X"06",X"1C",X"EA",X"07",X"0C",X"4B",X"27",X"60",X"AC",X"EA",X"02",X"B6",
		X"CF",X"F4",X"06",X"1C",X"EA",X"07",X"3E",X"7A",X"E1",X"01",X"3E",X"7A",X"C2",X"07",X"A4",X"B0",
		X"3C",X"6D",X"0F",X"F4",X"0F",X"ED",X"1D",X"D9",X"76",X"21",X"60",X"D9",X"19",X"00",X"4E",X"9B",
		X"14",X"08",X"D9",X"22",X"01",X"D9",X"21",X"06",X"F3",X"14",X"08",X"D9",X"22",X"02",X"D9",X"21",
		X"07",X"9B",X"98",X"08",X"4B",X"5F",X"60",X"19",X"B8",X"ED",X"30",X"4B",X"27",X"60",X"48",X"4B",
		X"28",X"60",X"57",X"4B",X"26",X"60",X"19",X"02",X"19",X"02",X"19",X"02",X"19",X"02",X"F4",X"02",
		X"7D",X"0D",X"2C",X"0F",X"F4",X"04",X"7D",X"0E",X"6A",X"6E",X"04",X"57",X"7A",X"6E",X"08",X"38",
		X"7A",X"6E",X"08",X"78",X"78",X"78",X"78",X"78",X"7A",X"6E",X"08",X"4B",X"28",X"60",X"76",X"97",
		X"61",X"AC",X"1C",X"57",X"08",X"B6",X"CF",X"F4",X"05",X"1C",X"88",X"08",X"4B",X"27",X"60",X"0C",
		X"AC",X"1C",X"66",X"08",X"B6",X"CF",X"F4",X"05",X"1C",X"88",X"08",X"0D",X"C0",X"69",X"A4",X"0A",
		X"3C",X"22",X"00",X"00",X"00",X"00",X"00",X"F4",X"63",X"9B",X"EA",X"0A",X"F4",X"59",X"2C",X"08",
		X"F4",X"62",X"E7",X"CC",X"09",X"9B",X"FE",X"09",X"7A",X"84",X"07",X"19",X"03",X"19",X"4A",X"A4",
		X"C7",X"1F",X"A4",X"8F",X"17",X"7A",X"F3",X"0A",X"76",X"21",X"60",X"19",X"03",X"19",X"4A",X"76",
		X"26",X"60",X"19",X"4A",X"76",X"00",X"60",X"19",X"54",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"25",
		X"05",X"DE",X"E1",X"61",X"A4",X"26",X"1F",X"F4",X"13",X"2C",X"02",X"25",X"12",X"97",X"5E",X"76",
		X"79",X"0C",X"B3",X"00",X"04",X"D6",X"FA",X"4B",X"65",X"60",X"F4",X"00",X"ED",X"06",X"D9",X"76",
		X"68",X"60",X"1A",X"04",X"D9",X"76",X"6B",X"60",X"D9",X"22",X"01",X"C8",X"99",X"D9",X"F8",X"01",
		X"D9",X"22",X"00",X"56",X"99",X"D9",X"F8",X"00",X"4B",X"65",X"60",X"F4",X"00",X"ED",X"05",X"76",
		X"C4",X"D2",X"1A",X"03",X"76",X"C3",X"D2",X"A4",X"06",X"1E",X"01",X"15",X"00",X"04",X"5E",X"72",
		X"5A",X"C6",X"76",X"F0",X"D1",X"F8",X"40",X"71",X"05",X"65",X"F4",X"06",X"2C",X"04",X"25",X"D9",
		X"1A",X"02",X"25",X"D8",X"76",X"10",X"D2",X"F8",X"40",X"71",X"05",X"B3",X"20",X"CB",X"A4",X"C7",
		X"1F",X"A4",X"8F",X"17",X"A4",X"5A",X"2D",X"DC",X"89",X"F3",X"76",X"F0",X"D1",X"71",X"FF",X"15",
		X"00",X"04",X"40",X"71",X"00",X"76",X"10",X"D2",X"71",X"FF",X"40",X"71",X"00",X"76",X"5F",X"60",
		X"19",X"FE",X"76",X"26",X"60",X"19",X"54",X"7A",X"84",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A4",X"2F",
		X"3F",X"A4",X"CD",X"3C",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"7A",X"62",X"06",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A4",X"E5",X"3F",X"A4",
		X"2B",X"3D",X"00",X"00",X"00",X"00",X"00",X"00",X"A4",X"BD",X"3D",X"66",X"26",X"CB",X"97",X"25",
		X"03",X"DE",X"3F",X"60",X"76",X"00",X"60",X"19",X"6E",X"A4",X"03",X"58",X"A4",X"89",X"49",X"01",
		X"DC",X"D3",X"3E",X"7A",X"84",X"07",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A4",X"E5",
		X"3F",X"66",X"76",X"0C",X"62",X"19",X"5A",X"76",X"01",X"60",X"19",X"5A",X"3E",X"A4",X"2B",X"3D",
		X"A4",X"BD",X"3D",X"F2",X"01",X"A4",X"2C",X"3C",X"7A",X"84",X"07",X"A4",X"C1",X"2A",X"76",X"00",
		X"60",X"19",X"FE",X"B5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A4",X"E5",X"3F",X"A4",X"2B",X"3D",
		X"A4",X"05",X"40",X"76",X"01",X"60",X"19",X"55",X"A4",X"64",X"2D",X"A4",X"CD",X"3C",X"66",X"76",
		X"5F",X"60",X"19",X"05",X"3E",X"F3",X"78",X"01",X"4B",X"65",X"60",X"F4",X"00",X"ED",X"13",X"4B",
		X"66",X"60",X"F4",X"00",X"ED",X"1F",X"4B",X"67",X"60",X"F4",X"00",X"9B",X"96",X"0B",X"25",X"01",
		X"1A",X"37",X"4B",X"67",X"60",X"F4",X"00",X"ED",X"0C",X"4B",X"66",X"60",X"F4",X"00",X"9B",X"96",
		X"0B",X"25",X"02",X"1A",X"24",X"4B",X"5F",X"60",X"19",X"04",X"7D",X"17",X"4B",X"65",X"60",X"F4",
		X"00",X"ED",X"09",X"4B",X"67",X"60",X"F4",X"00",X"ED",X"24",X"1A",X"07",X"4B",X"66",X"60",X"F4",
		X"00",X"ED",X"1B",X"7A",X"F7",X"21",X"FF",X"FF",X"FF",X"97",X"A4",X"99",X"3A",X"A4",X"F3",X"3C",
		X"00",X"00",X"00",X"01",X"A4",X"FC",X"2C",X"B3",X"80",X"A4",X"28",X"05",X"1A",X"09",X"A4",X"99",
		X"3A",X"A4",X"F3",X"3C",X"00",X"00",X"00",X"A4",X"74",X"2C",X"B3",X"80",X"A4",X"28",X"05",X"4B",
		X"65",X"60",X"8B",X"DE",X"65",X"60",X"A4",X"CD",X"3F",X"76",X"5F",X"60",X"19",X"0D",X"F3",X"0B",
		X"06",X"19",X"6E",X"7A",X"D5",X"04",X"A4",X"40",X"2B",X"B3",X"80",X"A4",X"28",X"05",X"76",X"1C",
		X"60",X"19",X"03",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"A4",X"BA",X"1A",X"A4",X"60",X"50",X"4B",
		X"5E",X"60",X"F4",X"00",X"7D",X"0A",X"76",X"02",X"90",X"19",X"86",X"7D",X"1D",X"7A",X"5F",X"03",
		X"76",X"02",X"90",X"19",X"86",X"7D",X"13",X"76",X"5F",X"60",X"19",X"03",X"B3",X"02",X"CB",X"B3",
		X"B4",X"A4",X"28",X"05",X"DC",X"89",X"F7",X"7A",X"1B",X"01",X"25",X"09",X"DE",X"5E",X"60",X"7A",
		X"5F",X"03",X"01",X"01",X"01",X"02",X"01",X"03",X"01",X"04",X"01",X"05",X"02",X"01",X"02",X"03",
		X"03",X"01",X"03",X"02",X"04",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"CA",X"D0",X"D0",X"D0",X"D6",X"D0",X"5A",X"D1",X"1A",X"D2",X"DA",X"D2",X"0A",X"D1",
		X"46",X"D1",X"4C",X"D1",X"D0",X"D1",X"12",X"D2",X"C6",X"D2",X"D4",X"D2",X"16",X"D3",X"4A",X"D3",
		X"50",X"D3",X"56",X"D3",X"06",X"D2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"10",X"15",X"20",X"25",X"30",X"35",X"40",
		X"45",X"50",X"55",X"60",X"65",X"70",X"75",X"80",X"85",X"90",X"95",X"18",X"30",X"60",X"48",X"78",
		X"90",X"A8",X"C0",X"12",X"15",X"15",X"16",X"15",X"12",X"17",X"12",X"17",X"18",X"1A",X"12",X"12",
		X"16",X"1B",X"15",X"16",X"17",X"5E",X"66",X"74",X"9A",X"63",X"72",X"8C",X"A2",X"62",X"70",X"88",
		X"A0",X"5B",X"64",X"74",X"94",X"59",X"64",X"74",X"90",X"5A",X"66",X"74",X"92",X"5C",X"64",X"74",
		X"96",X"5D",X"68",X"78",X"98",X"5C",X"6A",X"7C",X"96",X"5F",X"6C",X"80",X"9C",X"60",X"6E",X"84",
		X"9E",X"61",X"66",X"74",X"92",X"00",X"47",X"46",X"49",X"48",X"FF",X"4A",X"FF",X"00",X"41",X"39",
		X"00",X"40",X"42",X"43",X"00",X"44",X"45",X"01",X"39",X"01",X"35",X"36",X"37",X"01",X"FF",X"01",
		X"01",X"3D",X"01",X"40",X"3E",X"FF",X"01",X"3F",X"01",X"01",X"FC",X"06",X"F2",X"03",X"6D",X"06",
		X"C7",X"01",X"FC",X"03",X"6D",X"06",X"F2",X"06",X"C7",X"13",X"11",X"33",X"11",X"32",X"13",X"21",
		X"12",X"11",X"31",X"12",X"13",X"23",X"22",X"32",X"32",X"21",X"12",X"11",X"12",X"F5",X"D0",X"27",
		X"D1",X"2D",X"D1",X"39",X"D1",X"6F",X"D1",X"75",X"D1",X"A9",X"D1",X"AD",X"D1",X"B3",X"D1",X"B7",
		X"D1",X"69",X"D2",X"6D",X"D2",X"73",X"D2",X"77",X"D2",X"AF",X"D2",X"B5",X"D2",X"E7",X"D2",X"ED",
		X"D2",X"F9",X"D2",X"35",X"D3",X"32",X"3C",X"38",X"31",X"32",X"3B",X"38",X"33",X"33",X"3C",X"34",
		X"31",X"33",X"3B",X"34",X"33",X"20",X"01",X"13",X"12",X"20",X"11",X"33",X"33",X"12",X"10",X"FF",
		X"E5",X"5E",X"5B",X"59",X"5A",X"5C",X"5D",X"5C",X"5F",X"60",X"61",X"62",X"63",X"19",X"15",X"0A",
		X"22",X"0E",X"1B",X"FF",X"0C",X"11",X"0A",X"17",X"10",X"0E",X"02",X"02",X"02",X"01",X"01",X"01",
		X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"1C",
		X"21",X"2C",X"31",X"3E",X"43",X"49",X"56",X"5A",X"61",X"64",X"65",X"6A",X"6B",X"6C",X"6D",X"6E",
		X"6F",X"70",X"EC",X"EE",X"EE",X"EE",X"EE",X"06",X"FD",X"FF",X"FF",X"FF",X"FF",X"07",X"FD",X"FF",
		X"FF",X"FF",X"FF",X"07",X"FD",X"FF",X"FF",X"FF",X"FF",X"07",X"FD",X"FF",X"FF",X"FF",X"FF",X"07",
		X"FD",X"FF",X"FF",X"FF",X"FF",X"07",X"FD",X"FF",X"FF",X"FF",X"FF",X"07",X"FD",X"FF",X"FF",X"FF",
		X"FF",X"07",X"FD",X"FF",X"FF",X"FF",X"FF",X"07",X"FD",X"FF",X"FF",X"FF",X"FF",X"07",X"B9",X"BB",
		X"BB",X"BB",X"BB",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"02",X"03",X"05",X"03",X"06",X"09",X"15",X"08",X"16",X"24",X"40",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"33",X"FF",X"10",X"0A",X"16",X"0E",X"FF",X"18",X"1F",X"0E",
		X"1B",X"01",X"1C",X"1D",X"FF",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"02",X"17",X"0D",X"FF",X"19",
		X"15",X"0A",X"22",X"0E",X"1B",X"AE",X"AB",X"A7",X"AB",X"AE",X"A7",X"AB",X"00",X"01",X"02",X"03",
		X"00",X"03",X"03",X"03",X"04",X"00",X"04",X"04",X"04",X"04",X"00",X"04",X"05",X"05",X"05",X"00",
		X"06",X"06",X"06",X"07",X"90",X"24",X"00",X"00",X"02",X"04",X"01",X"03",X"05",X"06",X"08",X"05",
		X"07",X"09",X"0A",X"0B",X"08",X"0C",X"0D",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"12",X"12",X"12",X"15",X"15",X"15",X"18",X"18",
		X"18",X"18",X"18",X"20",X"20",X"20",X"20",X"20",X"12",X"12",X"15",X"15",X"18",X"18",X"18",X"18",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"08",X"08",X"04",X"04",X"04",X"02",X"02",
		X"02",X"04",X"04",X"04",X"02",X"02",X"02",X"04",X"04",X"08",X"08",X"08",X"08",X"08",X"01",X"01",
		X"01",X"08",X"08",X"08",X"01",X"01",X"01",X"08",X"08",X"08",X"08",X"08",X"04",X"04",X"02",X"02",
		X"02",X"04",X"04",X"08",X"08",X"04",X"04",X"08",X"08",X"04",X"04",X"02",X"02",X"01",X"01",X"01",
		X"01",X"01",X"02",X"02",X"01",X"01",X"01",X"08",X"08",X"08",X"01",X"01",X"01",X"01",X"01",X"02",
		X"02",X"04",X"04",X"04",X"02",X"02",X"02",X"04",X"04",X"04",X"02",X"02",X"02",X"02",X"02",X"02",
		X"02",X"02",X"01",X"01",X"08",X"08",X"08",X"01",X"01",X"02",X"02",X"01",X"01",X"02",X"02",X"01",
		X"01",X"08",X"08",X"08",X"08",X"04",X"04",X"08",X"08",X"08",X"08",X"01",X"01",X"08",X"08",X"04",
		X"04",X"02",X"02",X"02",X"04",X"04",X"04",X"02",X"02",X"02",X"04",X"04",X"04",X"02",X"02",X"02",
		X"04",X"04",X"04",X"02",X"02",X"01",X"01",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"04",X"04",
		X"04",X"04",X"04",X"08",X"FF",X"04",X"04",X"04",X"04",X"04",X"02",X"02",X"02",X"02",X"02",X"01",
		X"01",X"01",X"08",X"08",X"08",X"04",X"04",X"08",X"08",X"01",X"01",X"02",X"02",X"01",X"01",X"08",
		X"08",X"08",X"08",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"20",X"10",X"23",X"10",X"28",X"10",X"2D",X"10",X"30",X"10",X"33",X"10",X"36",X"10",X"3B",X"10",
		X"40",X"10",X"45",X"10",X"4A",X"10",X"4F",X"10",X"54",X"10",X"57",X"10",X"5C",X"10",X"5F",X"10",
		X"01",X"8B",X"10",X"02",X"C8",X"12",X"1D",X"13",X"02",X"88",X"12",X"A7",X"12",X"01",X"62",X"10",
		X"01",X"A7",X"10",X"01",X"A3",X"13",X"02",X"B9",X"10",X"00",X"11",X"02",X"47",X"11",X"56",X"11",
		X"02",X"DE",X"13",X"FF",X"13",X"02",X"65",X"11",X"76",X"11",X"02",X"0E",X"12",X"47",X"12",X"02",
		X"BC",X"11",X"E5",X"11",X"01",X"AC",X"10",X"02",X"87",X"11",X"16",X"14",X"01",X"9A",X"10",X"01",
		X"84",X"13",X"04",X"B0",X"05",X"C1",X"04",X"C2",X"04",X"C3",X"04",X"B1",X"05",X"C2",X"04",X"C3",
		X"04",X"C4",X"04",X"B2",X"05",X"C3",X"04",X"C4",X"04",X"C5",X"04",X"B3",X"05",X"C4",X"04",X"C5",
		X"04",X"C6",X"04",X"B4",X"05",X"C5",X"04",X"C6",X"04",X"C7",X"FF",X"30",X"C1",X"2F",X"C1",X"2D",
		X"C1",X"2B",X"C1",X"30",X"C1",X"30",X"C3",X"00",X"CF",X"FF",X"41",X"D0",X"00",X"EF",X"F1",X"F0",
		X"41",X"F0",X"41",X"F0",X"00",X"EF",X"FF",X"1C",X"F3",X"1F",X"F3",X"FF",X"1F",X"C0",X"23",X"C0",
		X"26",X"A0",X"23",X"A0",X"2B",X"80",X"00",X"AF",X"FF",X"2B",X"73",X"2A",X"A3",X"29",X"73",X"28",
		X"A3",X"26",X"93",X"24",X"C3",X"23",X"93",X"21",X"C3",X"1F",X"A3",X"00",X"CF",X"1F",X"C3",X"1E",
		X"93",X"1F",X"C3",X"21",X"93",X"1F",X"C3",X"1E",X"93",X"1F",X"C3",X"21",X"93",X"1F",X"C3",X"1E",
		X"93",X"1F",X"C3",X"28",X"A3",X"00",X"AF",X"28",X"63",X"1F",X"C3",X"1E",X"93",X"1F",X"C3",X"21",
		X"93",X"1F",X"C3",X"1E",X"93",X"1F",X"C3",X"21",X"83",X"23",X"83",X"24",X"53",X"00",X"EF",X"FF",
		X"13",X"72",X"12",X"A2",X"11",X"72",X"10",X"A2",X"0E",X"92",X"0C",X"C2",X"0B",X"92",X"09",X"C2",
		X"07",X"A2",X"00",X"CF",X"07",X"C2",X"06",X"92",X"07",X"C2",X"00",X"A2",X"00",X"AF",X"07",X"A2",
		X"00",X"AF",X"00",X"A2",X"00",X"AF",X"07",X"A2",X"00",X"AF",X"0C",X"A2",X"00",X"AF",X"0C",X"62",
		X"07",X"C2",X"06",X"92",X"07",X"C2",X"07",X"A2",X"00",X"AF",X"00",X"A2",X"00",X"AF",X"0C",X"82",
		X"0E",X"82",X"10",X"52",X"00",X"AF",X"FF",X"18",X"C1",X"1C",X"C1",X"1F",X"C1",X"24",X"C1",X"28",
		X"C1",X"2B",X"C1",X"30",X"C1",X"FF",X"13",X"C1",X"18",X"C1",X"1C",X"C1",X"1F",X"C1",X"24",X"C1",
		X"28",X"C1",X"2B",X"C1",X"FF",X"1B",X"D1",X"1D",X"D1",X"1F",X"D1",X"20",X"D1",X"22",X"D1",X"24",
		X"D1",X"26",X"D1",X"27",X"D1",X"FF",X"27",X"D1",X"26",X"D1",X"24",X"D1",X"22",X"D1",X"20",X"D1",
		X"1F",X"D1",X"1D",X"D1",X"1B",X"D1",X"FF",X"24",X"B2",X"26",X"B2",X"28",X"A2",X"00",X"CF",X"2B",
		X"A2",X"00",X"CF",X"2B",X"A2",X"00",X"CF",X"2D",X"A2",X"00",X"CF",X"2B",X"A2",X"00",X"CF",X"28",
		X"A2",X"00",X"CF",X"24",X"82",X"26",X"A2",X"28",X"A2",X"00",X"CF",X"28",X"A2",X"00",X"CF",X"26",
		X"A2",X"00",X"CF",X"26",X"A2",X"00",X"CF",X"24",X"92",X"00",X"CF",X"FF",X"28",X"83",X"2B",X"A3",
		X"28",X"A3",X"00",X"AF",X"26",X"A3",X"23",X"83",X"26",X"A3",X"23",X"A3",X"00",X"AF",X"1F",X"A3",
		X"21",X"83",X"1F",X"A3",X"1C",X"A3",X"00",X"8F",X"1C",X"73",X"0E",X"A3",X"00",X"AF",X"0E",X"A3",
		X"10",X"73",X"00",X"AF",X"FF",X"24",X"85",X"28",X"A5",X"24",X"A5",X"00",X"AF",X"23",X"A5",X"1F",
		X"85",X"23",X"A5",X"1F",X"A5",X"00",X"AF",X"1C",X"A5",X"1E",X"85",X"1C",X"A5",X"18",X"A5",X"00",
		X"8F",X"18",X"75",X"0B",X"A5",X"00",X"AF",X"0B",X"A5",X"0C",X"75",X"00",X"AF",X"FF",X"21",X"A2",
		X"23",X"C2",X"24",X"A2",X"00",X"AF",X"24",X"A2",X"00",X"AF",X"1F",X"A2",X"00",X"AF",X"1F",X"A2",
		X"00",X"AF",X"1C",X"A2",X"00",X"AF",X"1C",X"A2",X"00",X"AF",X"1A",X"82",X"18",X"92",X"1A",X"C2",
		X"1C",X"A2",X"1F",X"82",X"21",X"A2",X"1F",X"92",X"1C",X"C2",X"18",X"92",X"1A",X"C2",X"1C",X"82",
		X"1A",X"82",X"18",X"72",X"00",X"AF",X"FF",X"00",X"CF",X"00",X"AF",X"0C",X"A3",X"00",X"AF",X"13",
		X"A3",X"00",X"AF",X"0C",X"A3",X"00",X"AF",X"13",X"A3",X"00",X"AF",X"0C",X"A3",X"00",X"AF",X"13",
		X"A3",X"00",X"AF",X"13",X"A3",X"00",X"AF",X"0E",X"A3",X"00",X"AF",X"0C",X"A3",X"00",X"AF",X"13",
		X"A3",X"00",X"AF",X"0C",X"A3",X"00",X"AF",X"13",X"A3",X"00",X"AF",X"13",X"A3",X"00",X"AF",X"0E",
		X"A3",X"00",X"AF",X"0C",X"73",X"00",X"AF",X"FF",X"00",X"BF",X"30",X"C1",X"2F",X"C1",X"2D",X"C1",
		X"2B",X"C1",X"30",X"C1",X"2F",X"C1",X"2D",X"C1",X"2B",X"C1",X"30",X"C1",X"2F",X"C1",X"2D",X"C1",
		X"2B",X"C1",X"30",X"C1",X"30",X"C3",X"FF",X"00",X"BF",X"0C",X"C1",X"0B",X"C1",X"09",X"C1",X"07",
		X"C1",X"18",X"C1",X"17",X"C1",X"15",X"C1",X"13",X"C1",X"24",X"C1",X"23",X"C1",X"21",X"C1",X"1F",
		X"C1",X"24",X"C1",X"24",X"C3",X"00",X"AF",X"FF",X"1F",X"A3",X"21",X"93",X"22",X"C3",X"00",X"8F",
		X"23",X"A3",X"00",X"AF",X"1F",X"A3",X"00",X"AF",X"00",X"8F",X"23",X"83",X"00",X"AF",X"1F",X"A3",
		X"00",X"AF",X"1F",X"A3",X"21",X"93",X"23",X"C3",X"00",X"8F",X"24",X"A3",X"00",X"AF",X"1F",X"A3",
		X"00",X"7F",X"24",X"83",X"00",X"AF",X"1F",X"A3",X"00",X"AF",X"1F",X"A3",X"21",X"93",X"22",X"C3",
		X"00",X"8F",X"23",X"A3",X"00",X"AF",X"1F",X"A3",X"00",X"7F",X"23",X"83",X"00",X"AF",X"1F",X"A3",
		X"00",X"AF",X"1F",X"A3",X"21",X"93",X"23",X"C3",X"24",X"53",X"00",X"AF",X"FF",X"00",X"7F",X"0B",
		X"A4",X"00",X"AF",X"13",X"A4",X"00",X"AF",X"0B",X"A4",X"00",X"AF",X"13",X"A4",X"00",X"AF",X"0B",
		X"A4",X"00",X"AF",X"13",X"A4",X"00",X"AF",X"13",X"A4",X"00",X"AF",X"13",X"A4",X"00",X"AF",X"0C",
		X"A4",X"00",X"AF",X"13",X"A4",X"00",X"AF",X"0C",X"A4",X"00",X"AF",X"13",X"A4",X"00",X"AF",X"0C",
		X"A4",X"00",X"AF",X"13",X"A4",X"00",X"AF",X"0C",X"A4",X"00",X"AF",X"13",X"A4",X"00",X"AF",X"0B",
		X"A4",X"00",X"AF",X"13",X"A4",X"00",X"AF",X"0B",X"A4",X"00",X"AF",X"13",X"A4",X"00",X"AF",X"0B",
		X"A4",X"00",X"AF",X"13",X"A4",X"00",X"AF",X"10",X"A4",X"00",X"AF",X"13",X"A4",X"00",X"AF",X"0C",
		X"54",X"00",X"AF",X"FF",X"2D",X"E2",X"2A",X"E2",X"27",X"E2",X"24",X"E2",X"21",X"E2",X"1E",X"E2",
		X"1B",X"E2",X"18",X"E2",X"15",X"E2",X"12",X"E2",X"0F",X"E2",X"0C",X"E2",X"09",X"E2",X"06",X"E2",
		X"03",X"E2",X"FF",X"03",X"96",X"04",X"A5",X"05",X"B4",X"06",X"C3",X"07",X"D2",X"08",X"E1",X"03",
		X"96",X"04",X"A5",X"05",X"B4",X"06",X"C3",X"07",X"D2",X"08",X"E1",X"03",X"96",X"04",X"A5",X"05",
		X"B4",X"06",X"C3",X"07",X"D2",X"08",X"E1",X"03",X"96",X"04",X"A5",X"05",X"B4",X"06",X"C3",X"07",
		X"D2",X"08",X"E1",X"08",X"F4",X"07",X"F6",X"06",X"F8",X"05",X"FA",X"00",X"EF",X"FF",X"14",X"E0",
		X"15",X"E0",X"16",X"E1",X"17",X"E1",X"18",X"E2",X"19",X"E2",X"1A",X"E3",X"1B",X"E3",X"1C",X"E4",
		X"1D",X"E4",X"1E",X"E5",X"1F",X"E5",X"20",X"E6",X"21",X"E6",X"22",X"E7",X"00",X"EF",X"FF",X"81",
		X"E1",X"81",X"E1",X"81",X"E2",X"81",X"E3",X"81",X"E4",X"81",X"E5",X"81",X"E6",X"81",X"E7",X"81",
		X"E8",X"81",X"A9",X"00",X"EF",X"FF",X"1C",X"B2",X"1D",X"B2",X"1F",X"A2",X"00",X"CF",X"1C",X"A2",
		X"00",X"CF",X"1F",X"A2",X"00",X"CF",X"1C",X"A2",X"00",X"CF",X"1F",X"A2",X"00",X"CF",X"1C",X"A2",
		X"00",X"CF",X"1F",X"A2",X"00",X"CF",X"1C",X"A2",X"00",X"CF",X"1F",X"A2",X"00",X"CF",X"1F",X"A2",
		X"00",X"CF",X"1D",X"A2",X"00",X"CF",X"1D",X"A2",X"00",X"CF",X"18",X"96",X"13",X"96",X"0C",X"76",
		X"00",X"CF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"CB",X"72",X"25",X"01",X"23",X"7D",X"05",X"19",X"99",X"7A",X"36",X"17",X"DC",X"B5",
		X"26",X"97",X"65",X"5E",X"57",X"19",X"99",X"6B",X"D9",X"76",X"04",X"60",X"57",X"CE",X"00",X"D9",
		X"40",X"01",X"D3",X"B5",X"B5",X"76",X"00",X"70",X"B3",X"04",X"D4",X"00",X"CB",X"B3",X"FF",X"4B",
		X"01",X"90",X"19",X"F8",X"ED",X"F9",X"08",X"C0",X"89",X"F5",X"DC",X"89",X"EF",X"B5",X"25",X"9F",
		X"DE",X"00",X"B0",X"DE",X"00",X"C0",X"25",X"BF",X"DE",X"00",X"B0",X"DE",X"00",X"C0",X"25",X"DF",
		X"DE",X"00",X"B0",X"DE",X"00",X"C0",X"25",X"FF",X"DE",X"00",X"B0",X"DE",X"00",X"C0",X"B5",X"76",
		X"5F",X"60",X"19",X"05",X"9B",X"A1",X"17",X"76",X"00",X"60",X"EE",X"F8",X"C0",X"F8",X"C0",X"F8",
		X"B5",X"D9",X"66",X"76",X"00",X"60",X"22",X"6D",X"FF",X"F3",X"E5",X"17",X"C0",X"22",X"6D",X"FF",
		X"F3",X"D0",X"17",X"C0",X"22",X"6D",X"FF",X"9B",X"BF",X"18",X"B3",X"10",X"19",X"3D",X"1C",X"C4",
		X"17",X"A4",X"FA",X"17",X"14",X"32",X"65",X"F4",X"18",X"9B",X"BF",X"18",X"32",X"7A",X"BC",X"17",
		X"B3",X"08",X"19",X"3D",X"1C",X"DA",X"17",X"A4",X"FA",X"17",X"14",X"32",X"65",X"F4",X"10",X"7D",
		X"D2",X"32",X"7A",X"D2",X"17",X"B3",X"00",X"19",X"3D",X"1C",X"EF",X"17",X"A4",X"FA",X"17",X"14",
		X"32",X"65",X"F4",X"08",X"7D",X"B6",X"32",X"7A",X"E7",X"17",X"CB",X"97",X"66",X"76",X"00",X"10",
		X"19",X"ED",X"AE",X"B3",X"00",X"D6",X"3C",X"C0",X"FA",X"A5",X"E4",X"3C",X"C0",X"04",X"65",X"6D",
		X"FF",X"9B",X"AF",X"18",X"C2",X"69",X"C0",X"0D",X"C0",X"D9",X"76",X"03",X"60",X"7B",X"6D",X"C0",
		X"9B",X"46",X"18",X"D9",X"22",X"00",X"19",X"F8",X"ED",X"0C",X"B6",X"2F",X"16",X"60",X"D9",X"19",
		X"00",X"F6",X"23",X"7A",X"0D",X"18",X"23",X"19",X"B8",X"ED",X"D2",X"B6",X"2F",X"19",X"60",X"D9",
		X"19",X"00",X"FE",X"7A",X"0D",X"18",X"D9",X"22",X"00",X"19",X"72",X"F3",X"5A",X"18",X"B6",X"2F",
		X"04",X"60",X"D9",X"19",X"00",X"C6",X"23",X"7A",X"0D",X"18",X"19",X"04",X"F3",X"6B",X"18",X"B6",
		X"2F",X"07",X"60",X"D9",X"19",X"00",X"CE",X"23",X"7A",X"0D",X"18",X"19",X"48",X"F3",X"7C",X"18",
		X"B6",X"2F",X"0A",X"60",X"D9",X"19",X"00",X"D6",X"23",X"7A",X"0D",X"18",X"19",X"57",X"F3",X"8D",
		X"18",X"B6",X"2F",X"0D",X"60",X"D9",X"19",X"00",X"DE",X"23",X"7A",X"0D",X"18",X"19",X"E9",X"F3",
		X"9E",X"18",X"B6",X"2F",X"10",X"60",X"D9",X"19",X"00",X"E6",X"23",X"7A",X"0D",X"18",X"23",X"19",
		X"EB",X"F3",X"0D",X"18",X"B6",X"2F",X"13",X"60",X"D9",X"19",X"00",X"EE",X"7A",X"0D",X"18",X"3E",
		X"01",X"DC",X"32",X"65",X"6D",X"07",X"5C",X"A4",X"32",X"17",X"8B",X"CD",X"F8",X"32",X"B5",X"4B",
		X"03",X"60",X"B3",X"06",X"D9",X"76",X"04",X"60",X"19",X"02",X"E7",X"DA",X"18",X"D9",X"C0",X"D9",
		X"C0",X"D9",X"C0",X"23",X"9B",X"CF",X"19",X"7A",X"C8",X"18",X"32",X"D9",X"22",X"02",X"F4",X"00",
		X"7D",X"07",X"D9",X"9E",X"02",X"32",X"7A",X"CD",X"18",X"D9",X"24",X"00",X"D9",X"05",X"01",X"22",
		X"F4",X"FF",X"F3",X"3E",X"19",X"25",X"06",X"49",X"F4",X"03",X"2C",X"14",X"6E",X"03",X"19",X"99",
		X"19",X"99",X"19",X"99",X"19",X"99",X"19",X"99",X"FE",X"9F",X"DE",X"00",X"C0",X"7A",X"1F",X"19",
		X"19",X"99",X"19",X"99",X"19",X"99",X"19",X"99",X"19",X"99",X"FE",X"9F",X"DE",X"00",X"B0",X"25",
		X"06",X"49",X"48",X"F2",X"01",X"1D",X"F4",X"00",X"7D",X"06",X"2A",X"19",X"C0",X"7A",X"25",X"19",
		X"6A",X"8B",X"57",X"4B",X"03",X"60",X"8C",X"DE",X"03",X"60",X"32",X"7A",X"CD",X"18",X"25",X"06",
		X"49",X"F4",X"03",X"30",X"9A",X"19",X"6E",X"03",X"19",X"99",X"19",X"99",X"19",X"99",X"19",X"99",
		X"19",X"99",X"FE",X"80",X"04",X"E2",X"76",X"07",X"1B",X"22",X"6D",X"3F",X"19",X"99",X"57",X"CE",
		X"00",X"E2",X"40",X"E2",X"22",X"00",X"8F",X"DE",X"00",X"C0",X"E2",X"22",X"01",X"DE",X"00",X"C0",
		X"C0",X"25",X"00",X"B6",X"E9",X"8F",X"19",X"79",X"DE",X"00",X"C0",X"25",X"00",X"B6",X"EB",X"E2",
		X"76",X"F7",X"1A",X"C0",X"D9",X"1F",X"00",X"D9",X"C1",X"01",X"57",X"CE",X"00",X"E2",X"40",X"E2",
		X"22",X"00",X"5E",X"D9",X"F8",X"02",X"32",X"7A",X"CD",X"18",X"19",X"99",X"19",X"99",X"19",X"99",
		X"19",X"99",X"19",X"99",X"FE",X"80",X"04",X"E2",X"76",X"07",X"1B",X"22",X"6D",X"3F",X"19",X"99",
		X"57",X"CE",X"00",X"E2",X"40",X"E2",X"22",X"00",X"8F",X"DE",X"00",X"B0",X"E2",X"22",X"01",X"DE",
		X"00",X"B0",X"C0",X"EE",X"B6",X"E9",X"8F",X"19",X"79",X"DE",X"00",X"B0",X"7A",X"7B",X"19",X"19",
		X"02",X"2C",X"0D",X"D9",X"C0",X"D9",X"C0",X"D9",X"C0",X"19",X"02",X"2C",X"72",X"7A",X"B7",X"1A",
		X"32",X"D9",X"22",X"02",X"F4",X"00",X"7D",X"07",X"D9",X"9E",X"02",X"32",X"7A",X"D3",X"19",X"D9",
		X"24",X"00",X"D9",X"05",X"01",X"22",X"F4",X"FF",X"ED",X"11",X"25",X"FF",X"DE",X"00",X"B0",X"4B",
		X"03",X"60",X"6D",X"BF",X"DE",X"03",X"60",X"32",X"7A",X"D3",X"19",X"B3",X"00",X"19",X"02",X"19",
		X"89",X"19",X"02",X"19",X"02",X"19",X"02",X"19",X"02",X"19",X"02",X"5E",X"19",X"ED",X"19",X"ED",
		X"B2",X"FE",X"E0",X"DE",X"00",X"B0",X"C0",X"25",X"00",X"B6",X"E9",X"FE",X"F0",X"DE",X"00",X"B0",
		X"25",X"00",X"B6",X"EB",X"E2",X"76",X"F7",X"1A",X"C0",X"D9",X"1F",X"00",X"D9",X"C1",X"01",X"57",
		X"CE",X"00",X"E2",X"40",X"E2",X"22",X"00",X"5E",X"D9",X"F8",X"02",X"32",X"7A",X"D3",X"19",X"D9",
		X"22",X"02",X"F4",X"00",X"7D",X"06",X"D9",X"9E",X"02",X"7A",X"B7",X"1A",X"D9",X"24",X"00",X"D9",
		X"05",X"01",X"22",X"F4",X"FF",X"ED",X"10",X"25",X"FF",X"DE",X"00",X"C0",X"4B",X"03",X"60",X"6D",
		X"7F",X"DE",X"03",X"60",X"7A",X"B7",X"1A",X"B3",X"00",X"19",X"02",X"19",X"89",X"19",X"02",X"19",
		X"02",X"19",X"02",X"19",X"02",X"19",X"02",X"5E",X"19",X"ED",X"19",X"ED",X"B2",X"FE",X"E0",X"DE",
		X"00",X"C0",X"C0",X"25",X"00",X"B6",X"E9",X"FE",X"F0",X"DE",X"00",X"C0",X"25",X"00",X"B6",X"EB",
		X"E2",X"76",X"F7",X"1A",X"C0",X"D9",X"1F",X"00",X"D9",X"C1",X"01",X"57",X"CE",X"00",X"E2",X"40",
		X"E2",X"22",X"00",X"5E",X"D9",X"F8",X"02",X"D9",X"3E",X"B5",X"66",X"97",X"CB",X"76",X"80",X"D0",
		X"25",X"FF",X"D4",X"18",X"00",X"B3",X"20",X"F8",X"C0",X"89",X"FC",X"00",X"9A",X"F3",X"C4",X"1A",
		X"DC",X"01",X"3E",X"B5",X"25",X"00",X"B3",X"80",X"76",X"00",X"D0",X"F8",X"C0",X"89",X"FC",X"D4",
		X"00",X"B3",X"18",X"F8",X"15",X"20",X"00",X"40",X"89",X"F9",X"77",X"9A",X"F3",X"F6",X"1A",X"77",
		X"76",X"9F",X"D0",X"7A",X"E1",X"1A",X"B5",X"FF",X"C0",X"80",X"60",X"40",X"30",X"20",X"18",X"10",
		X"0C",X"08",X"06",X"04",X"03",X"02",X"01",X"08",X"3F",X"0F",X"3B",X"09",X"38",X"06",X"35",X"06",
		X"32",X"0A",X"2F",X"0E",X"2C",X"06",X"2A",X"00",X"28",X"0C",X"25",X"0A",X"23",X"0A",X"21",X"0C",
		X"1F",X"0F",X"1D",X"04",X"1C",X"0B",X"1A",X"03",X"19",X"0D",X"17",X"07",X"16",X"03",X"15",X"00",
		X"14",X"0E",X"12",X"0D",X"11",X"0D",X"10",X"0E",X"0F",X"00",X"0F",X"02",X"0E",X"06",X"0D",X"0A",
		X"0C",X"0E",X"0B",X"04",X"0B",X"0A",X"0A",X"00",X"0A",X"07",X"09",X"0F",X"08",X"07",X"08",X"0F",
		X"07",X"08",X"07",X"01",X"07",X"0B",X"06",X"05",X"06",X"0F",X"05",X"0A",X"05",X"05",X"05",X"00",
		X"05",X"0B",X"04",X"07",X"04",X"03",X"04",X"0F",X"03",X"0C",X"03",X"09",X"03",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"C1",X"15",X"19",X"17",X"B5",X"94",X"D4",X"00",X"CB",X"B3",X"00",X"A4",X"FC",X"1B",X"DC",
		X"89",X"02",X"1A",X"04",X"77",X"CB",X"1A",X"F2",X"00",X"00",X"00",X"B5",X"D9",X"76",X"55",X"0C",
		X"CE",X"00",X"65",X"F4",X"02",X"ED",X"02",X"F2",X"02",X"C2",X"19",X"99",X"19",X"99",X"26",X"CE",
		X"00",X"57",X"D9",X"40",X"D3",X"D9",X"69",X"00",X"CB",X"D9",X"3C",X"03",X"19",X"2C",X"19",X"2C",
		X"19",X"2C",X"19",X"2C",X"D9",X"24",X"01",X"D9",X"05",X"02",X"07",X"26",X"15",X"20",X"00",X"40",
		X"D3",X"89",X"F7",X"19",X"90",X"ED",X"15",X"78",X"D9",X"24",X"01",X"D9",X"05",X"02",X"C0",X"D9",
		X"3C",X"03",X"19",X"2C",X"19",X"2C",X"19",X"2C",X"19",X"2C",X"1A",X"DE",X"DC",X"65",X"F4",X"00",
		X"ED",X"17",X"14",X"CB",X"F7",X"20",X"00",X"D9",X"24",X"01",X"D9",X"05",X"02",X"D6",X"D9",X"22",
		X"03",X"6D",X"0F",X"72",X"F2",X"03",X"7A",X"2A",X"1C",X"B5",X"F7",X"00",X"00",X"76",X"9E",X"D0",
		X"25",X"4B",X"F8",X"D9",X"76",X"52",X"0C",X"D9",X"D6",X"D9",X"3C",X"00",X"A4",X"9B",X"1C",X"77",
		X"C2",X"F4",X"03",X"ED",X"EB",X"76",X"9D",X"D0",X"D9",X"76",X"61",X"0C",X"B3",X"18",X"15",X"20",
		X"00",X"D9",X"22",X"00",X"F8",X"D9",X"C0",X"40",X"89",X"F7",X"B5",X"5C",X"15",X"20",X"00",X"40",
		X"F8",X"40",X"89",X"FC",X"B5",X"C0",X"19",X"22",X"7D",X"FC",X"19",X"22",X"ED",X"FC",X"66",X"A4",
		X"3A",X"03",X"A4",X"8F",X"17",X"3E",X"19",X"22",X"7D",X"FC",X"B5",X"CB",X"72",X"25",X"01",X"89",
		X"02",X"DC",X"B5",X"06",X"1A",X"F7",X"B5",X"00",X"4B",X"62",X"60",X"F4",X"00",X"7D",X"04",X"F2",
		X"06",X"1A",X"02",X"F2",X"05",X"D4",X"00",X"B3",X"0C",X"76",X"1C",X"D6",X"07",X"A4",X"24",X"1D",
		X"14",X"25",X"17",X"33",X"ED",X"0A",X"77",X"25",X"04",X"67",X"ED",X"02",X"D4",X"00",X"B3",X"00",
		X"25",X"00",X"67",X"ED",X"05",X"25",X"0C",X"33",X"7D",X"1E",X"4B",X"60",X"60",X"67",X"ED",X"15",
		X"4B",X"61",X"60",X"33",X"ED",X"0F",X"37",X"63",X"60",X"78",X"4B",X"62",X"60",X"F4",X"00",X"7D",
		X"03",X"38",X"1A",X"01",X"7C",X"7A",X"DC",X"1C",X"EE",X"DD",X"ED",X"07",X"4B",X"62",X"60",X"8B",
		X"DE",X"62",X"60",X"B5",X"26",X"19",X"42",X"7D",X"0A",X"19",X"39",X"7D",X"03",X"C0",X"1A",X"10",
		X"0C",X"1A",X"0D",X"19",X"39",X"7D",X"05",X"15",X"E0",X"FF",X"1A",X"03",X"15",X"20",X"00",X"40",
		X"D3",X"B5",X"25",X"52",X"D4",X"00",X"76",X"9C",X"D0",X"32",X"25",X"4E",X"B3",X"16",X"F8",X"A4",
		X"24",X"1D",X"32",X"F8",X"A4",X"24",X"1D",X"89",X"FA",X"F4",X"55",X"7D",X"06",X"5C",X"32",X"5C",
		X"77",X"1A",X"E9",X"B5",X"15",X"20",X"00",X"76",X"A3",X"D4",X"25",X"06",X"B3",X"0C",X"F8",X"66",
		X"C0",X"F8",X"3E",X"40",X"89",X"F8",X"B5",X"15",X"20",X"00",X"4B",X"65",X"60",X"F4",X"00",X"7D",
		X"05",X"4B",X"67",X"60",X"1A",X"03",X"4B",X"66",X"60",X"F4",X"07",X"2C",X"02",X"25",X"06",X"72",
		X"EE",X"32",X"25",X"06",X"49",X"04",X"CB",X"76",X"A3",X"D0",X"25",X"E1",X"DE",X"C8",X"61",X"EE",
		X"33",X"4B",X"C8",X"61",X"7D",X"08",X"F8",X"5C",X"40",X"F8",X"5E",X"40",X"89",X"F8",X"25",X"FF",
		X"42",X"19",X"ED",X"DE",X"C8",X"61",X"EE",X"33",X"4B",X"C8",X"61",X"7D",X"04",X"F8",X"40",X"89",
		X"FC",X"32",X"F4",X"FF",X"7D",X"0A",X"8B",X"32",X"76",X"A4",X"D0",X"25",X"E3",X"DC",X"1A",X"CC",
		X"B5",X"EE",X"A4",X"4C",X"1E",X"15",X"20",X"00",X"4B",X"5F",X"60",X"19",X"04",X"7D",X"13",X"76",
		X"43",X"D2",X"71",X"02",X"40",X"71",X"1E",X"40",X"7A",X"31",X"49",X"D9",X"76",X"6B",X"60",X"A4",
		X"06",X"1E",X"76",X"44",X"D2",X"71",X"01",X"40",X"71",X"1E",X"40",X"7A",X"3A",X"49",X"D9",X"76",
		X"68",X"60",X"A4",X"06",X"1E",X"B5",X"26",X"CB",X"66",X"B3",X"03",X"76",X"DA",X"61",X"66",X"D9",
		X"22",X"00",X"04",X"19",X"02",X"19",X"02",X"19",X"02",X"19",X"02",X"F8",X"C0",X"C2",X"6D",X"0F",
		X"F8",X"D9",X"C0",X"C0",X"89",X"E9",X"3E",X"B3",X"05",X"EE",X"21",X"ED",X"05",X"71",X"FF",X"C0",
		X"89",X"F8",X"3E",X"D9",X"66",X"D9",X"76",X"DA",X"61",X"15",X"20",X"00",X"B3",X"06",X"D9",X"22",
		X"00",X"F8",X"D9",X"C0",X"40",X"89",X"F7",X"D9",X"3E",X"DC",X"D3",X"B5",X"97",X"CB",X"66",X"F4",
		X"00",X"ED",X"14",X"25",X"03",X"76",X"44",X"D6",X"B3",X"0A",X"A4",X"7D",X"1E",X"76",X"43",X"D6",
		X"B3",X"0A",X"A4",X"7D",X"1E",X"1A",X"12",X"4B",X"65",X"60",X"F4",X"00",X"ED",X"07",X"76",X"44",
		X"D6",X"25",X"00",X"1A",X"EB",X"25",X"00",X"1A",X"E4",X"3E",X"DC",X"01",X"B5",X"CB",X"26",X"66",
		X"15",X"20",X"00",X"F8",X"40",X"89",X"FC",X"3E",X"D3",X"DC",X"B5",X"76",X"E2",X"D4",X"25",X"06",
		X"B3",X"08",X"A4",X"7D",X"1E",X"76",X"E2",X"D0",X"71",X"11",X"15",X"20",X"00",X"40",X"71",X"12",
		X"40",X"71",X"2A",X"40",X"A4",X"24",X"5F",X"A4",X"BD",X"25",X"B5",X"8B",X"FF",X"BC",X"3F",X"77",
		X"1A",X"17",X"FF",X"FF",X"FF",X"FF",X"FF",X"B3",X"09",X"76",X"80",X"D3",X"D9",X"76",X"AB",X"1E",
		X"CB",X"B3",X"03",X"D9",X"22",X"00",X"F8",X"C0",X"D9",X"C0",X"89",X"F7",X"DC",X"89",X"ED",X"B3",
		X"09",X"76",X"73",X"60",X"71",X"01",X"C0",X"71",X"00",X"C0",X"71",X"00",X"C0",X"89",X"F5",X"B5",
		X"76",X"E1",X"D0",X"15",X"20",X"00",X"71",X"1B",X"40",X"71",X"18",X"40",X"71",X"1E",X"40",X"71",
		X"17",X"7A",X"1D",X"5F",X"76",X"A1",X"D1",X"15",X"20",X"00",X"A4",X"26",X"1F",X"F4",X"00",X"7D",
		X"24",X"F4",X"64",X"2C",X"08",X"71",X"09",X"40",X"71",X"09",X"7A",X"25",X"1F",X"B3",X"00",X"D4",
		X"0A",X"67",X"2C",X"04",X"82",X"14",X"1A",X"F9",X"32",X"EE",X"33",X"7D",X"03",X"A3",X"1A",X"02",
		X"71",X"FF",X"40",X"32",X"F8",X"B5",X"4B",X"65",X"60",X"19",X"04",X"7D",X"05",X"4B",X"6F",X"60",
		X"1A",X"03",X"4B",X"6E",X"60",X"B5",X"4B",X"02",X"90",X"19",X"B8",X"7D",X"04",X"25",X"03",X"1A",
		X"02",X"25",X"05",X"B5",X"A4",X"26",X"1F",X"F4",X"00",X"ED",X"04",X"71",X"FF",X"1A",X"2F",X"5E",
		X"F4",X"12",X"2C",X"02",X"25",X"11",X"CE",X"00",X"57",X"E2",X"76",X"79",X"0C",X"E2",X"40",X"15",
		X"20",X"00",X"E2",X"22",X"00",X"04",X"6D",X"F0",X"7D",X"0A",X"19",X"02",X"19",X"02",X"19",X"02",
		X"19",X"02",X"F8",X"40",X"C2",X"6D",X"0F",X"F8",X"40",X"71",X"00",X"40",X"71",X"00",X"B5",X"D9",
		X"66",X"A4",X"26",X"1F",X"F4",X"00",X"7D",X"07",X"5E",X"F4",X"12",X"2C",X"02",X"25",X"11",X"D9",
		X"76",X"93",X"0C",X"04",X"B3",X"00",X"D9",X"D6",X"D9",X"3C",X"00",X"D4",X"00",X"19",X"99",X"19",
		X"99",X"C8",X"D9",X"3E",X"B5",X"D9",X"22",X"01",X"F4",X"07",X"1C",X"AF",X"1F",X"25",X"07",X"6E",
		X"07",X"57",X"19",X"73",X"19",X"73",X"19",X"73",X"19",X"73",X"6D",X"0F",X"32",X"6A",X"F4",X"0B",
		X"E7",X"C5",X"1F",X"F2",X"0B",X"32",X"B5",X"D9",X"66",X"A4",X"7D",X"44",X"A4",X"5A",X"2D",X"76",
		X"01",X"90",X"19",X"22",X"9B",X"D2",X"1F",X"76",X"59",X"60",X"D1",X"22",X"76",X"5A",X"60",X"6D",
		X"03",X"ED",X"01",X"D1",X"A4",X"3A",X"03",X"76",X"4E",X"60",X"EE",X"B3",X"0B",X"F8",X"C0",X"89",
		X"FC",X"D9",X"76",X"1C",X"60",X"D9",X"22",X"00",X"6D",X"03",X"F3",X"0C",X"20",X"14",X"25",X"0A");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
