library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_cpu2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_cpu2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"33",X"9B",X"03",X"21",X"15",X"05",X"00",X"D9",X"40",X"7A",X"F5",X"1F",X"76",X"5F",X"60",X"19",
		X"FA",X"7D",X"20",X"76",X"02",X"90",X"19",X"24",X"7D",X"19",X"04",X"4B",X"65",X"60",X"F4",X"00",
		X"C2",X"7D",X"10",X"D9",X"FA",X"02",X"25",X"FE",X"82",X"04",X"D9",X"0D",X"01",X"25",X"AE",X"DA",
		X"7A",X"39",X"20",X"D9",X"22",X"01",X"D9",X"FA",X"02",X"D9",X"0D",X"00",X"19",X"4B",X"19",X"4B",
		X"19",X"4B",X"19",X"4B",X"A4",X"40",X"22",X"26",X"CE",X"00",X"E2",X"76",X"4E",X"60",X"E2",X"40",
		X"97",X"E2",X"22",X"00",X"E2",X"D1",X"00",X"CB",X"8D",X"14",X"E2",X"76",X"80",X"70",X"15",X"40",
		X"00",X"E2",X"40",X"89",X"FC",X"19",X"99",X"19",X"99",X"57",X"E2",X"40",X"DC",X"C2",X"6E",X"07",
		X"E2",X"F8",X"03",X"01",X"6D",X"0F",X"D3",X"F2",X"00",X"19",X"29",X"ED",X"06",X"19",X"90",X"7D",
		X"06",X"19",X"79",X"7C",X"7A",X"8D",X"20",X"19",X"E8",X"ED",X"02",X"19",X"68",X"76",X"5F",X"60",
		X"19",X"FA",X"7D",X"2A",X"76",X"02",X"90",X"19",X"24",X"7D",X"23",X"DE",X"C8",X"61",X"4B",X"65",
		X"60",X"F4",X"00",X"4B",X"C8",X"61",X"7D",X"16",X"19",X"E9",X"ED",X"05",X"19",X"79",X"7A",X"B3",
		X"20",X"19",X"0A",X"19",X"EB",X"ED",X"05",X"19",X"68",X"7A",X"BE",X"20",X"19",X"EE",X"FE",X"C0",
		X"E2",X"F8",X"00",X"D9",X"22",X"03",X"D9",X"19",X"04",X"66",X"ED",X"2B",X"F4",X"D8",X"EA",X"27",
		X"32",X"EE",X"4C",X"ED",X"06",X"32",X"5A",X"0C",X"7A",X"DC",X"20",X"32",X"32",X"4B",X"5A",X"60",
		X"6D",X"03",X"19",X"72",X"7D",X"05",X"CE",X"04",X"7A",X"F1",X"20",X"F4",X"02",X"ED",X"07",X"CE",
		X"08",X"32",X"EC",X"7A",X"F7",X"20",X"32",X"E2",X"F8",X"01",X"D9",X"22",X"04",X"E2",X"F8",X"02",
		X"7A",X"FD",X"1F",X"76",X"C0",X"70",X"B3",X"0B",X"D9",X"76",X"4E",X"60",X"D9",X"22",X"00",X"66",
		X"19",X"99",X"19",X"99",X"57",X"CE",X"00",X"40",X"91",X"66",X"D3",X"6A",X"D3",X"26",X"A2",X"F4",
		X"20",X"EA",X"0D",X"E2",X"3E",X"E2",X"66",X"15",X"20",X"00",X"E2",X"40",X"EE",X"E2",X"F8",X"00",
		X"15",X"40",X"00",X"D9",X"C0",X"3E",X"40",X"89",X"D3",X"76",X"01",X"90",X"19",X"22",X"F3",X"3C",
		X"21",X"D9",X"3E",X"B5",X"25",X"00",X"B3",X"16",X"76",X"A6",X"D4",X"15",X"20",X"00",X"CB",X"B3",
		X"16",X"66",X"F8",X"C0",X"89",X"FC",X"3E",X"DC",X"40",X"89",X"F3",X"B5",X"B5",X"FF",X"FF",X"FF",
		X"26",X"CB",X"97",X"A4",X"CC",X"56",X"4B",X"0F",X"62",X"F4",X"AA",X"7D",X"09",X"01",X"DC",X"D3",
		X"76",X"2B",X"60",X"7A",X"BA",X"07",X"25",X"00",X"DE",X"0F",X"62",X"A4",X"84",X"57",X"2C",X"06",
		X"01",X"DC",X"D3",X"7A",X"53",X"22",X"76",X"D1",X"57",X"3C",X"D4",X"00",X"C0",X"22",X"CB",X"66",
		X"76",X"F9",X"D4",X"A4",X"23",X"56",X"22",X"3E",X"DC",X"6D",X"0F",X"F4",X"03",X"ED",X"01",X"77",
		X"89",X"EA",X"19",X"4F",X"4B",X"3B",X"62",X"67",X"EA",X"C3",X"F4",X"0B",X"EA",X"BF",X"76",X"3B",
		X"62",X"D1",X"C0",X"D1",X"4B",X"3B",X"62",X"76",X"BE",X"D0",X"F7",X"40",X"00",X"D6",X"5E",X"ED",
		X"FC",X"15",X"00",X"04",X"66",X"71",X"53",X"0C",X"71",X"E7",X"0C",X"71",X"E6",X"3E",X"40",X"71",
		X"02",X"0C",X"71",X"02",X"0C",X"71",X"02",X"25",X"D7",X"16",X"ED",X"18",X"25",X"7C",X"3A",X"ED",
		X"13",X"71",X"02",X"C0",X"71",X"02",X"C0",X"71",X"02",X"76",X"7C",X"D3",X"71",X"4F",X"C0",X"71",
		X"4F",X"C0",X"71",X"4E",X"7A",X"6D",X"21",X"A4",X"FD",X"21",X"7A",X"DC",X"04",X"25",X"00",X"DE",
		X"C9",X"61",X"15",X"54",X"54",X"25",X"02",X"B3",X"0B",X"76",X"BE",X"D0",X"A4",X"D1",X"5D",X"15",
		X"FF",X"FF",X"25",X"02",X"B3",X"0B",X"76",X"BD",X"D0",X"A4",X"D1",X"5D",X"15",X"E5",X"E5",X"25",
		X"02",X"B3",X"0B",X"76",X"BC",X"D0",X"A4",X"D1",X"5D",X"76",X"7C",X"D3",X"71",X"4F",X"C0",X"71",
		X"4F",X"C0",X"71",X"4E",X"76",X"7C",X"D7",X"71",X"02",X"C0",X"71",X"02",X"C0",X"71",X"02",X"B5",
		X"97",X"1D",X"F4",X"02",X"ED",X"09",X"4B",X"4B",X"62",X"F4",X"00",X"ED",X"02",X"CE",X"08",X"01",
		X"7A",X"A8",X"1F",X"B3",X"80",X"A4",X"73",X"22",X"76",X"01",X"60",X"19",X"6E",X"A4",X"2F",X"3F",
		X"B3",X"30",X"A4",X"73",X"22",X"00",X"00",X"A4",X"64",X"4B",X"76",X"F8",X"0E",X"37",X"D8",X"61",
		X"7A",X"A0",X"22",X"CB",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"DC",X"89",X"F6",X"B5",X"66",X"76",
		X"5F",X"60",X"19",X"05",X"7D",X"06",X"3E",X"71",X"02",X"7A",X"FB",X"35",X"3E",X"F4",X"01",X"ED",
		X"05",X"71",X"02",X"7A",X"FB",X"35",X"F4",X"05",X"1C",X"F1",X"35",X"71",X"03",X"7A",X"FB",X"35",
		X"A4",X"FD",X"21",X"7A",X"5E",X"09",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"66",X"CB",X"B3",X"FF",X"CB",X"B3",X"FF",X"CB",X"B3",X"FF",X"00",
		X"89",X"FD",X"DC",X"89",X"F7",X"DC",X"89",X"F1",X"DC",X"3E",X"B5",X"66",X"CB",X"66",X"F4",X"04",
		X"2C",X"10",X"19",X"72",X"7D",X"06",X"E2",X"76",X"F0",X"0C",X"1A",X"52",X"E2",X"76",X"E7",X"0C",
		X"1A",X"4C",X"D4",X"00",X"19",X"72",X"7D",X"24",X"15",X"E1",X"FF",X"40",X"32",X"22",X"F4",X"E5",
		X"ED",X"02",X"19",X"DC",X"15",X"3E",X"00",X"40",X"22",X"F4",X"E5",X"ED",X"02",X"19",X"70",X"97",
		X"C2",X"DE",X"8E",X"60",X"01",X"32",X"E2",X"76",X"DE",X"0C",X"1A",X"22",X"15",X"21",X"00",X"40",
		X"32",X"22",X"F4",X"E5",X"ED",X"02",X"19",X"B5",X"15",X"BE",X"FF",X"40",X"22",X"F4",X"E5",X"ED",
		X"02",X"19",X"D3",X"97",X"C2",X"DE",X"8E",X"60",X"01",X"32",X"E2",X"76",X"D5",X"0C",X"A4",X"0F",
		X"24",X"3E",X"D4",X"00",X"32",X"19",X"4B",X"19",X"9D",X"1C",X"DF",X"23",X"C2",X"F4",X"00",X"ED",
		X"05",X"A4",X"D9",X"24",X"1A",X"79",X"F4",X"04",X"ED",X"05",X"A4",X"8B",X"24",X"1A",X"70",X"A4",
		X"23",X"24",X"26",X"E2",X"66",X"CE",X"00",X"5E",X"F4",X"04",X"2C",X"01",X"5E",X"57",X"E2",X"40",
		X"E2",X"22",X"00",X"E2",X"3E",X"D3",X"F4",X"01",X"ED",X"40",X"66",X"76",X"8E",X"60",X"C2",X"F4",
		X"03",X"ED",X"06",X"19",X"FA",X"7D",X"18",X"1A",X"1A",X"EA",X"06",X"19",X"3C",X"7D",X"10",X"1A",
		X"12",X"F4",X"08",X"ED",X"06",X"19",X"0D",X"7D",X"06",X"1A",X"08",X"19",X"69",X"ED",X"04",X"25",
		X"FF",X"1A",X"14",X"25",X"E5",X"97",X"25",X"02",X"D9",X"66",X"26",X"15",X"00",X"04",X"D9",X"40",
		X"D9",X"F8",X"00",X"D3",X"D9",X"3E",X"01",X"3E",X"1A",X"12",X"97",X"25",X"05",X"D9",X"66",X"26",
		X"15",X"00",X"04",X"D9",X"40",X"D9",X"F8",X"00",X"D3",X"D9",X"3E",X"01",X"D9",X"F8",X"00",X"C2",
		X"F4",X"0A",X"7D",X"05",X"77",X"32",X"7A",X"54",X"23",X"32",X"F4",X"04",X"2C",X"0D",X"25",X"00",
		X"DE",X"8E",X"60",X"DE",X"90",X"60",X"DE",X"8F",X"60",X"1A",X"11",X"25",X"09",X"DE",X"8F",X"60",
		X"25",X"01",X"DE",X"90",X"60",X"66",X"76",X"00",X"60",X"19",X"5A",X"3E",X"DC",X"3E",X"B5",X"97",
		X"19",X"99",X"57",X"CE",X"00",X"D9",X"76",X"F9",X"0C",X"D9",X"40",X"D9",X"0D",X"00",X"D9",X"69",
		X"01",X"01",X"B5",X"26",X"66",X"D9",X"3E",X"F4",X"06",X"7D",X"3C",X"F4",X"02",X"ED",X"04",X"D9",
		X"C0",X"1A",X"34",X"EA",X"07",X"15",X"E1",X"FF",X"D9",X"40",X"1A",X"2B",X"F4",X"05",X"ED",X"05",
		X"15",X"E0",X"FF",X"1A",X"F3",X"EA",X"05",X"15",X"21",X"00",X"1A",X"EC",X"F4",X"08",X"ED",X"05",
		X"15",X"DF",X"FF",X"1A",X"E3",X"EA",X"05",X"15",X"20",X"00",X"1A",X"DC",X"F4",X"09",X"7D",X"05",
		X"15",X"1F",X"00",X"1A",X"D3",X"D9",X"0C",X"D3",X"B5",X"7A",X"A9",X"56",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"26",X"66",X"15",X"C0",X"FF",
		X"40",X"A4",X"69",X"24",X"F4",X"02",X"ED",X"0D",X"32",X"F4",X"04",X"2C",X"04",X"71",X"34",X"1A",
		X"34",X"71",X"33",X"1A",X"30",X"EA",X"0D",X"32",X"F4",X"04",X"2C",X"04",X"71",X"38",X"1A",X"25",
		X"71",X"FF",X"1A",X"21",X"32",X"F4",X"04",X"2C",X"0E",X"32",X"22",X"F4",X"3B",X"ED",X"04",X"71",
		X"3A",X"1A",X"13",X"71",X"34",X"1A",X"0F",X"32",X"22",X"F4",X"3A",X"ED",X"04",X"71",X"3B",X"1A",
		X"05",X"71",X"33",X"1A",X"01",X"32",X"3E",X"D3",X"B5",X"26",X"66",X"C0",X"C0",X"A4",X"69",X"24",
		X"F4",X"02",X"ED",X"0D",X"32",X"F4",X"04",X"2C",X"04",X"71",X"3B",X"1A",X"34",X"71",X"33",X"1A",
		X"30",X"EA",X"0D",X"32",X"F4",X"04",X"2C",X"04",X"71",X"3C",X"1A",X"25",X"71",X"FF",X"1A",X"21",
		X"32",X"F4",X"04",X"2C",X"0E",X"32",X"22",X"F4",X"34",X"ED",X"04",X"71",X"3A",X"1A",X"13",X"71",
		X"3B",X"1A",X"0F",X"32",X"22",X"F4",X"3A",X"ED",X"04",X"71",X"34",X"1A",X"05",X"71",X"33",X"1A",
		X"01",X"32",X"3E",X"D3",X"B5",X"A4",X"06",X"2B",X"A4",X"BA",X"1A",X"A4",X"55",X"17",X"A4",X"3E",
		X"25",X"A4",X"60",X"4C",X"A4",X"1D",X"27",X"A4",X"CB",X"27",X"A4",X"26",X"28",X"B5",X"B3",X"10",
		X"76",X"1E",X"D1",X"D9",X"76",X"D7",X"2E",X"D4",X"04",X"A4",X"B3",X"27",X"76",X"1C",X"D1",X"B3",
		X"01",X"66",X"65",X"F4",X"01",X"7D",X"08",X"D4",X"03",X"A4",X"B1",X"25",X"F8",X"1A",X"07",X"D4",
		X"00",X"A4",X"B1",X"25",X"71",X"1D",X"15",X"20",X"00",X"40",X"D9",X"76",X"CF",X"2E",X"F4",X"05",
		X"EA",X"08",X"5E",X"19",X"99",X"CE",X"00",X"57",X"1A",X"03",X"15",X"06",X"00",X"D9",X"40",X"A4",
		X"B1",X"25",X"D9",X"22",X"00",X"F8",X"D9",X"C0",X"26",X"15",X"20",X"00",X"40",X"D3",X"A4",X"B1",
		X"25",X"D9",X"22",X"00",X"F8",X"26",X"15",X"40",X"00",X"40",X"D3",X"A4",X"BD",X"25",X"3E",X"14",
		X"65",X"F4",X"0A",X"EA",X"0B",X"F4",X"02",X"ED",X"04",X"0C",X"0C",X"1A",X"A4",X"0C",X"1A",X"A1",
		X"B5",X"97",X"66",X"26",X"15",X"00",X"04",X"40",X"08",X"D3",X"3E",X"01",X"B5",X"CB",X"D9",X"76",
		X"80",X"D3",X"65",X"5E",X"72",X"7D",X"05",X"EE",X"5A",X"08",X"89",X"FC",X"57",X"CE",X"00",X"D9",
		X"40",X"B3",X"07",X"15",X"00",X"04",X"66",X"40",X"08",X"3E",X"D9",X"22",X"00",X"F8",X"26",X"15",
		X"20",X"00",X"40",X"D9",X"C0",X"D3",X"89",X"EE",X"B3",X"06",X"C2",X"66",X"40",X"A4",X"7D",X"1E",
		X"3E",X"DC",X"D9",X"76",X"73",X"60",X"65",X"CB",X"5E",X"72",X"19",X"99",X"17",X"DC",X"57",X"CE",
		X"00",X"D9",X"40",X"A4",X"06",X"1E",X"B5",X"B5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"97",X"66",X"F8",X"5C",X"66",X"40",X"F8",X"3E",X"0C",X"5C",
		X"F8",X"40",X"5C",X"F8",X"3E",X"01",X"B5",X"CB",X"B3",X"03",X"F8",X"5C",X"40",X"89",X"FB",X"DC",
		X"B5",X"CB",X"B3",X"03",X"F8",X"5E",X"0A",X"B6",X"29",X"89",X"F9",X"DC",X"B5",X"B3",X"09",X"76",
		X"8B",X"D1",X"D9",X"76",X"F1",X"2E",X"D4",X"03",X"00",X"00",X"00",X"B3",X"02",X"76",X"EA",X"D1",
		X"D9",X"76",X"FA",X"2E",X"D4",X"03",X"00",X"00",X"00",X"B3",X"0E",X"76",X"29",X"D1",X"D9",X"76",
		X"FC",X"2E",X"D4",X"03",X"A4",X"B3",X"27",X"B3",X"05",X"76",X"C7",X"D1",X"D9",X"76",X"0A",X"2F",
		X"D4",X"01",X"A4",X"B3",X"27",X"4B",X"02",X"90",X"19",X"F8",X"ED",X"33",X"B3",X"03",X"76",X"06",
		X"D1",X"D9",X"76",X"21",X"2F",X"D4",X"01",X"A4",X"B3",X"27",X"B3",X"0E",X"76",X"86",X"D1",X"D9",
		X"76",X"24",X"2F",X"A4",X"B3",X"27",X"15",X"00",X"04",X"76",X"C6",X"D0",X"D4",X"04",X"66",X"40",
		X"08",X"3E",X"71",X"01",X"76",X"66",X"D1",X"66",X"40",X"08",X"3E",X"71",X"02",X"1A",X"23",X"4B",
		X"5E",X"60",X"F4",X"01",X"ED",X"C6",X"15",X"00",X"04",X"76",X"C6",X"D0",X"D4",X"04",X"66",X"40",
		X"08",X"3E",X"71",X"01",X"B3",X"12",X"76",X"06",X"D1",X"D9",X"76",X"0F",X"2F",X"D4",X"01",X"A4",
		X"B3",X"27",X"B5",X"26",X"15",X"00",X"04",X"66",X"40",X"08",X"3E",X"D9",X"22",X"00",X"F8",X"26",
		X"15",X"20",X"00",X"40",X"D9",X"C0",X"D3",X"89",X"EE",X"D3",X"B5",X"97",X"CB",X"26",X"66",X"B3",
		X"09",X"76",X"82",X"D4",X"25",X"02",X"15",X"20",X"00",X"F8",X"C0",X"F8",X"40",X"F8",X"0C",X"F8",
		X"40",X"89",X"F6",X"1A",X"07",X"97",X"CB",X"26",X"66",X"15",X"20",X"00",X"4B",X"5E",X"60",X"72",
		X"25",X"09",X"33",X"1A",X"1C",X"EE",X"76",X"03",X"90",X"B6",X"EB",X"76",X"82",X"D0",X"F4",X"0F",
		X"ED",X"0B",X"D4",X"E9",X"C2",X"A4",X"16",X"28",X"40",X"89",X"F9",X"1A",X"04",X"D4",X"ED",X"1A",
		X"F3",X"3E",X"D3",X"DC",X"01",X"B5",X"26",X"15",X"20",X"00",X"F8",X"5E",X"C0",X"F8",X"5E",X"40",
		X"F8",X"5E",X"0C",X"F8",X"D3",X"B5",X"15",X"20",X"00",X"B3",X"08",X"76",X"81",X"D6",X"25",X"02",
		X"F8",X"40",X"89",X"FC",X"4B",X"02",X"90",X"19",X"F8",X"7D",X"1B",X"B3",X"06",X"D9",X"76",X"81",
		X"D2",X"76",X"E7",X"2E",X"A4",X"CF",X"29",X"76",X"61",X"D3",X"4B",X"5E",X"60",X"F4",X"09",X"2C",
		X"02",X"25",X"09",X"F8",X"1A",X"0C",X"B3",X"04",X"D9",X"76",X"01",X"D3",X"76",X"ED",X"2E",X"A4",
		X"CF",X"29",X"B5",X"B5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"66",X"A4",
		X"1C",X"29",X"A4",X"C1",X"2A",X"76",X"B3",X"D1",X"A4",X"E3",X"1E",X"A4",X"82",X"29",X"A4",X"A8",
		X"29",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3E",X"B5",X"76",X"B3",X"D5",X"25",
		X"05",X"B3",X"05",X"A4",X"74",X"29",X"76",X"D5",X"D5",X"25",X"01",X"23",X"A4",X"74",X"29",X"76",
		X"74",X"D5",X"25",X"04",X"B3",X"0A",X"A4",X"74",X"29",X"76",X"33",X"D5",X"25",X"00",X"B3",X"0F",
		X"00",X"00",X"00",X"76",X"10",X"D5",X"25",X"03",X"B3",X"10",X"A4",X"74",X"29",X"C0",X"A4",X"74",
		X"29",X"76",X"AD",X"D5",X"25",X"05",X"B3",X"06",X"A4",X"74",X"29",X"C0",X"A4",X"74",X"29",X"76",
		X"AA",X"D5",X"A4",X"74",X"29",X"C0",X"A4",X"74",X"29",X"76",X"10",X"D5",X"25",X"03",X"B3",X"10",
		X"A4",X"74",X"29",X"B5",X"CB",X"66",X"97",X"15",X"20",X"00",X"F8",X"40",X"89",X"FC",X"01",X"3E",
		X"DC",X"B5",X"76",X"D5",X"D1",X"71",X"FF",X"15",X"20",X"00",X"40",X"00",X"00",X"00",X"D9",X"76",
		X"21",X"60",X"D9",X"71",X"00",X"82",X"D9",X"71",X"01",X"58",X"D9",X"71",X"02",X"AE",X"A4",X"7F",
		X"1F",X"D9",X"F8",X"03",X"D9",X"A3",X"04",X"B5",X"A4",X"26",X"1F",X"B3",X"11",X"76",X"4A",X"2F",
		X"15",X"0F",X"00",X"5E",X"7D",X"03",X"40",X"89",X"FA",X"D9",X"76",X"33",X"D1",X"B3",X"0F",X"00",
		X"00",X"00",X"B3",X"10",X"D9",X"76",X"10",X"D1",X"76",X"50",X"30",X"A4",X"CF",X"29",X"B5",X"26",
		X"15",X"20",X"00",X"22",X"D9",X"F8",X"00",X"C0",X"D9",X"40",X"89",X"F7",X"D3",X"B5",X"A4",X"26",
		X"1F",X"76",X"B0",X"D2",X"F4",X"12",X"2C",X"07",X"B3",X"06",X"A4",X"32",X"2A",X"1A",X"42",X"F4",
		X"0A",X"2C",X"0D",X"B3",X"05",X"15",X"20",X"00",X"0A",X"B6",X"29",X"A4",X"32",X"2A",X"1A",X"31",
		X"F4",X"05",X"2C",X"0D",X"B3",X"04",X"15",X"40",X"00",X"0A",X"B6",X"29",X"A4",X"32",X"2A",X"1A",
		X"20",X"F4",X"02",X"2C",X"0D",X"B3",X"03",X"15",X"60",X"00",X"0A",X"B6",X"29",X"A4",X"32",X"2A",
		X"1A",X"0F",X"F4",X"01",X"2C",X"0B",X"B3",X"02",X"15",X"80",X"00",X"0A",X"B6",X"29",X"A4",X"32",
		X"2A",X"B5",X"15",X"20",X"00",X"71",X"63",X"C0",X"71",X"73",X"0A",X"B6",X"29",X"71",X"F0",X"0C",
		X"71",X"A3",X"0A",X"B6",X"29",X"89",X"EE",X"B5",X"76",X"4D",X"D2",X"E2",X"76",X"6F",X"60",X"B3",
		X"03",X"D9",X"76",X"AD",X"0C",X"E2",X"C0",X"E2",X"69",X"00",X"19",X"C0",X"19",X"C0",X"CE",X"00",
		X"D9",X"40",X"A4",X"68",X"2A",X"89",X"EA",X"B5",X"26",X"15",X"20",X"00",X"D9",X"22",X"00",X"F8",
		X"C0",X"D9",X"C0",X"D9",X"22",X"00",X"5C",X"F8",X"0A",X"B6",X"29",X"A4",X"91",X"2A",X"F8",X"0C",
		X"D9",X"C0",X"D9",X"C0",X"D9",X"22",X"00",X"5C",X"F8",X"15",X"20",X"00",X"0A",X"B6",X"29",X"D3",
		X"B5",X"CB",X"E2",X"22",X"00",X"B3",X"F1",X"F4",X"09",X"7D",X"08",X"6E",X"05",X"2C",X"04",X"5C",
		X"17",X"1A",X"01",X"65",X"DC",X"B5",X"76",X"4A",X"D2",X"B3",X"03",X"15",X"20",X"00",X"71",X"62",
		X"C0",X"71",X"71",X"0A",X"B6",X"29",X"71",X"EF",X"0C",X"71",X"A1",X"0A",X"B6",X"29",X"89",X"EE",
		X"B5",X"A4",X"FD",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"76",X"A6",X"D0",X"15",X"20",X"00",X"25",X"FF",X"D4",X"16",X"66",X"B3",
		X"16",X"F8",X"40",X"89",X"FC",X"3E",X"C0",X"9A",X"ED",X"F4",X"B5",X"66",X"26",X"15",X"00",X"04",
		X"40",X"71",X"00",X"D3",X"3E",X"B5",X"F7",X"FF",X"03",X"76",X"00",X"D4",X"EE",X"F8",X"C0",X"D0",
		X"65",X"8F",X"ED",X"F8",X"B5",X"76",X"0B",X"62",X"15",X"0C",X"00",X"B3",X"0A",X"71",X"00",X"C0",
		X"71",X"00",X"C0",X"71",X"00",X"C0",X"71",X"00",X"C0",X"71",X"00",X"40",X"89",X"EF",X"A4",X"C7",
		X"1F",X"7A",X"C1",X"54",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"66",X"76",X"AB",X"62",X"71",X"00",X"C0",X"71",X"00",X"C0",X"71",X"00",X"3E",X"7A",X"FC",X"2C",
		X"15",X"00",X"04",X"CB",X"FA",X"C0",X"3C",X"C0",X"66",X"CB",X"3E",X"40",X"F8",X"C0",X"F8",X"26",
		X"15",X"E0",X"FF",X"40",X"F8",X"0C",X"F8",X"D3",X"3E",X"DC",X"89",X"E7",X"B5",X"76",X"99",X"61",
		X"D1",X"22",X"97",X"76",X"A8",X"61",X"B3",X"06",X"6D",X"0F",X"F4",X"00",X"ED",X"07",X"25",X"02",
		X"A4",X"50",X"2B",X"1A",X"09",X"F4",X"08",X"ED",X"05",X"25",X"01",X"A4",X"50",X"2B",X"01",X"97",
		X"6D",X"07",X"76",X"A2",X"61",X"B3",X"03",X"F4",X"00",X"ED",X"05",X"A4",X"C6",X"2B",X"1A",X"07",
		X"F4",X"04",X"ED",X"03",X"A4",X"C6",X"2B",X"01",X"97",X"6D",X"1F",X"76",X"9C",X"61",X"B3",X"03",
		X"F4",X"00",X"ED",X"07",X"25",X"00",X"A4",X"50",X"2B",X"1A",X"09",X"F4",X"10",X"ED",X"05",X"25",
		X"03",X"A4",X"50",X"2B",X"01",X"B5",X"CB",X"FA",X"C0",X"3C",X"C0",X"66",X"CB",X"3E",X"15",X"E1",
		X"FF",X"40",X"22",X"15",X"20",X"00",X"F4",X"7F",X"ED",X"10",X"71",X"7B",X"0C",X"71",X"7A",X"40",
		X"71",X"5D",X"C0",X"71",X"78",X"3E",X"DC",X"89",X"DD",X"B5",X"F4",X"83",X"ED",X"0D",X"71",X"7F",
		X"0C",X"71",X"7E",X"40",X"71",X"5C",X"C0",X"71",X"7C",X"1A",X"EA",X"F4",X"77",X"ED",X"0D",X"71",
		X"83",X"0C",X"71",X"82",X"40",X"71",X"5B",X"C0",X"71",X"80",X"1A",X"D9",X"F4",X"7B",X"ED",X"0D",
		X"71",X"77",X"0C",X"71",X"9A",X"40",X"71",X"5E",X"C0",X"71",X"66",X"1A",X"C8",X"F4",X"79",X"ED",
		X"04",X"71",X"74",X"1A",X"ED",X"F4",X"7D",X"ED",X"04",X"71",X"79",X"1A",X"AF",X"F4",X"81",X"ED",
		X"04",X"71",X"7D",X"1A",X"BB",X"71",X"81",X"1A",X"C8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"1D",X"F4",X"00",X"7D",X"0C",X"F4",
		X"02",X"7D",X"0C",X"F4",X"03",X"ED",X"0A",X"71",X"3B",X"1A",X"06",X"71",X"34",X"1A",X"02",X"71",
		X"3A",X"CE",X"00",X"B5",X"A4",X"C1",X"2A",X"76",X"26",X"60",X"19",X"FA",X"7D",X"03",X"A4",X"A2",
		X"2C",X"76",X"50",X"D1",X"25",X"FF",X"B3",X"0D",X"A4",X"7D",X"1E",X"76",X"50",X"D5",X"25",X"06",
		X"B3",X"0D",X"A4",X"7D",X"1E",X"76",X"6D",X"0D",X"D9",X"76",X"50",X"D1",X"B3",X"0D",X"A4",X"CF",
		X"29",X"B5",X"EE",X"76",X"21",X"60",X"F8",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"76",X"2B",X"60",
		X"B3",X"07",X"15",X"05",X"00",X"EE",X"F8",X"26",X"A4",X"4F",X"2E",X"D3",X"40",X"89",X"F7",X"76",
		X"26",X"60",X"66",X"71",X"12",X"C0",X"A4",X"4F",X"2E",X"9E",X"22",X"F4",X"07",X"ED",X"F7",X"3E",
		X"71",X"22",X"C0",X"C0",X"A4",X"4F",X"2E",X"9E",X"22",X"F4",X"22",X"ED",X"F7",X"76",X"26",X"60",
		X"71",X"00",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"4B",X"65",X"60",X"F4",X"00",X"7D",X"05",X"76",
		X"67",X"60",X"1A",X"03",X"76",X"66",X"60",X"D1",X"A4",X"77",X"1D",X"B5",X"97",X"A4",X"C1",X"2A",
		X"76",X"71",X"D5",X"B3",X"0A",X"25",X"00",X"A4",X"7D",X"1E",X"0C",X"A4",X"7D",X"1E",X"0C",X"A4",
		X"7D",X"1E",X"01",X"F4",X"01",X"7D",X"10",X"EA",X"28",X"B3",X"09",X"D9",X"76",X"90",X"D1",X"76",
		X"68",X"0E",X"A4",X"CF",X"29",X"1A",X"32",X"B3",X"0A",X"D9",X"76",X"71",X"D1",X"76",X"71",X"0E",
		X"A4",X"CF",X"29",X"B3",X"09",X"D9",X"76",X"8F",X"D1",X"76",X"68",X"0E",X"A4",X"CF",X"29",X"1A",
		X"18",X"B3",X"0A",X"D9",X"76",X"71",X"D1",X"76",X"7B",X"0E",X"A4",X"CF",X"29",X"B3",X"09",X"D9",
		X"76",X"8F",X"D1",X"76",X"68",X"0E",X"A4",X"CF",X"29",X"B5",X"97",X"4B",X"02",X"90",X"19",X"E9",
		X"7D",X"F9",X"01",X"B5",X"76",X"26",X"60",X"71",X"82",X"B3",X"1E",X"25",X"48",X"C0",X"C0",X"C0",
		X"A4",X"4F",X"2E",X"F8",X"C0",X"71",X"10",X"0C",X"89",X"F6",X"B3",X"03",X"5A",X"04",X"D4",X"08",
		X"F8",X"A4",X"4F",X"2E",X"9A",X"ED",X"F9",X"89",X"F3",X"B3",X"04",X"25",X"58",X"D4",X"18",X"F8",
		X"C0",X"71",X"10",X"19",X"6D",X"0C",X"A4",X"4F",X"2E",X"9A",X"ED",X"F3",X"5A",X"04",X"89",X"ED",
		X"B3",X"1E",X"F8",X"A4",X"4F",X"2E",X"89",X"FA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"15",X"CE",X"2D",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D3",X"76",X"26",
		X"60",X"71",X"00",X"A4",X"2F",X"3F",X"B5",X"0C",X"B3",X"02",X"25",X"AF",X"D1",X"21",X"9B",X"12",
		X"2E",X"A4",X"4F",X"2E",X"89",X"F6",X"B3",X"04",X"25",X"AF",X"D1",X"21",X"9B",X"12",X"2E",X"C0",
		X"D1",X"25",X"D7",X"21",X"9B",X"12",X"2E",X"A4",X"4F",X"2E",X"0C",X"89",X"EB",X"C0",X"B3",X"04",
		X"D1",X"21",X"9B",X"12",X"2E",X"A4",X"4F",X"2E",X"89",X"F6",X"B3",X"05",X"A4",X"4F",X"2E",X"89",
		X"FB",X"B5",X"D3",X"B5",X"0C",X"B3",X"02",X"EE",X"9E",X"21",X"9B",X"4D",X"2E",X"A4",X"4F",X"2E",
		X"89",X"F6",X"B3",X"04",X"EE",X"9E",X"21",X"9B",X"4D",X"2E",X"C0",X"D1",X"25",X"D7",X"21",X"9B",
		X"4D",X"2E",X"A4",X"4F",X"2E",X"0C",X"89",X"EC",X"C0",X"B3",X"04",X"D1",X"21",X"9B",X"4D",X"2E",
		X"A4",X"4F",X"2E",X"89",X"F6",X"B3",X"05",X"A4",X"4F",X"2E",X"89",X"FB",X"B5",X"D3",X"B5",X"97",
		X"66",X"CB",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"DC",X"3E",X"01",X"B5",X"76",X"A4",X"0E",X"A4",
		X"26",X"1F",X"19",X"72",X"ED",X"01",X"C0",X"4B",X"B9",X"61",X"21",X"E7",X"9E",X"2E",X"4B",X"65",
		X"60",X"F4",X"00",X"7D",X"0C",X"4B",X"02",X"90",X"19",X"EB",X"7D",X"05",X"4B",X"01",X"90",X"1A",
		X"03",X"4B",X"00",X"90",X"F4",X"00",X"9B",X"9E",X"2E",X"4B",X"98",X"61",X"76",X"C4",X"61",X"B3",
		X"04",X"19",X"02",X"EA",X"02",X"19",X"75",X"F8",X"C0",X"89",X"F6",X"7A",X"CB",X"2E",X"76",X"C4",
		X"61",X"B3",X"04",X"B6",X"57",X"6D",X"0F",X"19",X"02",X"5C",X"F4",X"03",X"2C",X"0D",X"F4",X"05",
		X"2C",X"0E",X"F4",X"07",X"2C",X"0F",X"25",X"08",X"7A",X"C7",X"2E",X"25",X"01",X"7A",X"C7",X"2E",
		X"25",X"02",X"7A",X"C7",X"2E",X"25",X"04",X"F8",X"C0",X"89",X"D8",X"A4",X"31",X"30",X"B5",X"18",
		X"19",X"17",X"0D",X"1B",X"0D",X"1D",X"11",X"1D",X"18",X"0D",X"0A",X"22",X"2E",X"1C",X"FF",X"11",
		X"12",X"2A",X"1C",X"0C",X"18",X"1B",X"0E",X"0C",X"1B",X"0E",X"0D",X"12",X"1D",X"0F",X"1B",X"0E",
		X"0E",X"19",X"1B",X"0E",X"1C",X"0E",X"17",X"1D",X"0E",X"0D",X"0B",X"22",X"2F",X"FF",X"01",X"09",
		X"08",X"03",X"FF",X"0F",X"0A",X"15",X"0C",X"18",X"17",X"FF",X"19",X"1E",X"1C",X"11",X"FF",X"19",
		X"15",X"0A",X"22",X"0E",X"1B",X"FF",X"0B",X"1E",X"1D",X"1D",X"18",X"17",X"FF",X"18",X"17",X"15",
		X"22",X"18",X"1B",X"FF",X"FF",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"FF",X"0B",X"1E",X"1D",X"1D",
		X"18",X"17",X"C0",X"AB",X"C1",X"A8",X"A8",X"C1",X"B9",X"C3",X"B2",X"C2",X"AB",X"C0",X"BD",X"C4",
		X"C5",X"AF",X"C2",X"B2",X"B9",X"C3",X"BD",X"C4",X"A8",X"C1",X"D9",X"66",X"76",X"0C",X"62",X"19",
		X"3C",X"7D",X"13",X"D9",X"76",X"2B",X"60",X"15",X"05",X"00",X"B3",X"04",X"D9",X"19",X"00",X"4E",
		X"ED",X"0A",X"D9",X"40",X"89",X"F6",X"19",X"03",X"B3",X"1E",X"1A",X"09",X"19",X"FA",X"74",X"AE",
		X"2F",X"ED",X"F3",X"B3",X"48",X"D9",X"3E",X"CB",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"A4",X"5A",
		X"2D",X"76",X"0C",X"62",X"19",X"3C",X"74",X"8D",X"2F",X"DC",X"89",X"EB",X"B5",X"3E",X"DC",X"CB",
		X"66",X"65",X"F4",X"01",X"ED",X"28",X"76",X"0C",X"62",X"5C",X"F8",X"4B",X"C3",X"61",X"0C",X"F8",
		X"25",X"10",X"DE",X"C3",X"61",X"A4",X"AE",X"2F",X"25",X"48",X"D4",X"03",X"1A",X"22",X"97",X"EE",
		X"DE",X"60",X"60",X"5C",X"DE",X"99",X"61",X"25",X"0D",X"DE",X"61",X"60",X"01",X"B5",X"BC",X"84",
		X"BC",X"84",X"BC",X"84",X"6D",X"0F",X"31",X"72",X"25",X"68",X"5A",X"04",X"89",X"FC",X"D4",X"1C",
		X"D9",X"66",X"D9",X"76",X"2B",X"60",X"15",X"05",X"00",X"B3",X"04",X"D9",X"19",X"00",X"4E",X"7D",
		X"06",X"D9",X"F8",X"03",X"D9",X"08",X"04",X"D9",X"40",X"89",X"F0",X"D9",X"3E",X"B5",X"FF",X"FF",
		X"4B",X"0C",X"62",X"19",X"57",X"ED",X"06",X"A4",X"3F",X"3E",X"7A",X"F8",X"3D",X"66",X"76",X"27",
		X"60",X"3C",X"C0",X"22",X"76",X"0C",X"62",X"19",X"12",X"3E",X"7A",X"FB",X"3D",X"D9",X"66",X"D9",
		X"76",X"2B",X"60",X"76",X"0C",X"62",X"15",X"05",X"00",X"B3",X"04",X"25",X"48",X"D9",X"19",X"00",
		X"4E",X"7D",X"05",X"D9",X"21",X"03",X"7D",X"06",X"D9",X"40",X"89",X"F1",X"19",X"AC",X"D9",X"3E",
		X"B5",X"4B",X"0C",X"62",X"19",X"04",X"E6",X"D8",X"46",X"B5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0C",X"11",X"0A",X"17",X"10",X"0E",X"FF",X"1D",X"18",X"FF",X"20",X"11",X"12",X"1D",X"0E",X"28",
		X"FF",X"C2",X"D9",X"76",X"2B",X"60",X"19",X"99",X"19",X"99",X"C8",X"CE",X"00",X"57",X"D9",X"40",
		X"D9",X"71",X"00",X"82",X"D9",X"71",X"01",X"58",X"D9",X"71",X"02",X"86",X"D9",X"71",X"03",X"18",
		X"D9",X"71",X"04",X"03",X"B5",X"FF",X"FF",X"97",X"66",X"A4",X"26",X"1F",X"5E",X"6D",X"07",X"76",
		X"8B",X"0C",X"CE",X"00",X"57",X"40",X"FA",X"76",X"A0",X"30",X"40",X"3C",X"3E",X"01",X"C2",X"B5",
		X"94",X"94",X"94",X"94",X"94",X"94",X"94",X"94",X"76",X"0C",X"62",X"19",X"FA",X"7D",X"04",X"19",
		X"4A",X"19",X"6E",X"76",X"2B",X"60",X"B5",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A4",
		X"A9",X"34",X"72",X"25",X"75",X"49",X"DE",X"A9",X"60",X"B5",X"B3",X"03",X"4B",X"65",X"60",X"F4",
		X"00",X"7D",X"05",X"76",X"A6",X"60",X"1A",X"03",X"76",X"A3",X"60",X"71",X"95",X"C0",X"71",X"6A",
		X"C0",X"71",X"0A",X"B5",X"4B",X"65",X"60",X"F4",X"00",X"7D",X"05",X"4B",X"A0",X"60",X"1A",X"03",
		X"4B",X"9D",X"60",X"B3",X"07",X"76",X"BD",X"D4",X"CE",X"03",X"F2",X"07",X"3D",X"2C",X"03",X"00",
		X"1A",X"01",X"91",X"26",X"15",X"20",X"00",X"40",X"D3",X"89",X"F1",X"B5",X"4B",X"65",X"60",X"F4",
		X"00",X"7D",X"05",X"4B",X"A1",X"60",X"1A",X"03",X"4B",X"9E",X"60",X"B3",X"05",X"76",X"DD",X"D5",
		X"CE",X"03",X"F2",X"06",X"3D",X"2C",X"03",X"07",X"1A",X"01",X"91",X"26",X"15",X"20",X"00",X"40",
		X"D3",X"89",X"F1",X"B5",X"76",X"9F",X"60",X"4B",X"65",X"60",X"F4",X"00",X"7D",X"03",X"76",X"A2",
		X"60",X"EE",X"F8",X"B5",X"4B",X"65",X"60",X"F4",X"00",X"7D",X"05",X"4B",X"A2",X"60",X"1A",X"03",
		X"4B",X"9F",X"60",X"76",X"BD",X"D6",X"15",X"20",X"00",X"B3",X"03",X"D4",X"05",X"F4",X"00",X"ED",
		X"0D",X"A3",X"40",X"A3",X"40",X"A3",X"40",X"A3",X"40",X"A3",X"40",X"A3",X"1A",X"13",X"08",X"40",
		X"08",X"F4",X"01",X"7D",X"EF",X"40",X"08",X"40",X"08",X"F4",X"02",X"7D",X"EB",X"40",X"08",X"40",
		X"08",X"B5",X"A4",X"63",X"33",X"A4",X"3D",X"3F",X"B3",X"0A",X"CE",X"00",X"E2",X"76",X"91",X"60",
		X"E2",X"66",X"E2",X"22",X"01",X"A4",X"C5",X"32",X"E2",X"C0",X"E2",X"C0",X"E2",X"C0",X"E2",X"C0",
		X"78",X"25",X"03",X"DD",X"ED",X"EC",X"A4",X"A9",X"34",X"E2",X"3E",X"B3",X"0B",X"CE",X"00",X"32",
		X"E2",X"22",X"02",X"A4",X"C5",X"32",X"E2",X"C0",X"E2",X"C0",X"E2",X"C0",X"E2",X"C0",X"78",X"32",
		X"5E",X"7D",X"0E",X"32",X"1D",X"F4",X"03",X"ED",X"E7",X"E2",X"76",X"92",X"60",X"CE",X"00",X"1A",
		X"DF",X"CE",X"00",X"E2",X"76",X"70",X"60",X"B6",X"57",X"06",X"19",X"18",X"06",X"6D",X"03",X"50",
		X"CE",X"00",X"F4",X"01",X"1A",X"32",X"2C",X"10",X"F4",X"03",X"9B",X"68",X"7A",X"30",X"78",X"32",
		X"F4",X"0D",X"30",X"A7",X"32",X"7A",X"88",X"32",X"E2",X"3C",X"00",X"4B",X"91",X"60",X"A4",X"C5",
		X"32",X"78",X"E2",X"3C",X"01",X"4B",X"95",X"60",X"A4",X"C5",X"32",X"78",X"E2",X"3C",X"02",X"4B",
		X"99",X"60",X"A4",X"C5",X"32",X"7A",X"C4",X"32",X"E2",X"3C",X"00",X"4B",X"91",X"60",X"A4",X"C5",
		X"32",X"78",X"E2",X"3C",X"02",X"4B",X"95",X"60",X"A4",X"C5",X"32",X"78",X"E2",X"3C",X"01",X"4B",
		X"99",X"60",X"A4",X"C5",X"32",X"7A",X"C4",X"32",X"E2",X"3C",X"01",X"4B",X"91",X"60",X"A4",X"C5",
		X"32",X"78",X"E2",X"3C",X"00",X"4B",X"95",X"60",X"A4",X"C5",X"32",X"78",X"E2",X"3C",X"02",X"4B",
		X"99",X"60",X"A4",X"C5",X"32",X"7A",X"C4",X"32",X"E2",X"3C",X"01",X"4B",X"91",X"60",X"A4",X"C5",
		X"32",X"78",X"E2",X"3C",X"02",X"4B",X"95",X"60",X"A4",X"C5",X"32",X"78",X"E2",X"3C",X"00",X"4B",
		X"99",X"60",X"A4",X"C5",X"32",X"7A",X"C4",X"32",X"E2",X"3C",X"02",X"4B",X"91",X"60",X"A4",X"C5",
		X"32",X"78",X"E2",X"3C",X"00",X"4B",X"95",X"60",X"A4",X"C5",X"32",X"78",X"E2",X"3C",X"01",X"4B",
		X"99",X"60",X"A4",X"C5",X"32",X"1A",X"1D",X"E2",X"3C",X"02",X"4B",X"91",X"60",X"A4",X"C5",X"32",
		X"78",X"E2",X"3C",X"01",X"4B",X"95",X"60",X"A4",X"C5",X"32",X"78",X"E2",X"3C",X"00",X"4B",X"99",
		X"60",X"A4",X"C5",X"32",X"B5",X"97",X"A4",X"79",X"3A",X"A4",X"44",X"34",X"01",X"97",X"CB",X"04",
		X"1D",X"A4",X"3B",X"33",X"DC",X"65",X"1A",X"01",X"97",X"CB",X"B3",X"03",X"F4",X"0A",X"ED",X"06",
		X"D9",X"76",X"A5",X"0C",X"1A",X"0A",X"F4",X"0B",X"ED",X"09",X"B3",X"01",X"D9",X"76",X"A9",X"0C",
		X"26",X"1A",X"0E",X"D9",X"76",X"AD",X"0C",X"26",X"19",X"99",X"19",X"99",X"CE",X"00",X"57",X"00",
		X"00",X"D9",X"22",X"00",X"F8",X"15",X"00",X"04",X"66",X"40",X"A3",X"3E",X"D9",X"22",X"01",X"C0",
		X"00",X"00",X"00",X"00",X"00",X"F8",X"66",X"40",X"A3",X"3E",X"26",X"15",X"E0",X"FF",X"40",X"D3",
		X"D9",X"22",X"02",X"C8",X"F8",X"66",X"40",X"A3",X"3E",X"0C",X"D9",X"22",X"03",X"19",X"42",X"7D",
		X"01",X"5C",X"F8",X"66",X"40",X"A3",X"3E",X"D3",X"DC",X"01",X"B5",X"D9",X"66",X"CB",X"F4",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"02",X"0C",X"1A",X"03",X"00",X"00",
		X"00",X"B3",X"00",X"19",X"76",X"D6",X"66",X"D9",X"3E",X"D9",X"24",X"00",X"D9",X"05",X"01",X"DC",
		X"D9",X"3E",X"B5",X"B3",X"0C",X"7A",X"B5",X"33",X"66",X"D9",X"3E",X"B6",X"57",X"04",X"BC",X"C3",
		X"6D",X"0F",X"19",X"76",X"19",X"76",X"54",X"00",X"A4",X"82",X"33",X"2C",X"EE",X"F8",X"C0",X"89",
		X"EA",X"B5",X"66",X"CB",X"47",X"76",X"91",X"60",X"21",X"7D",X"10",X"C0",X"97",X"92",X"5E",X"67",
		X"7D",X"03",X"01",X"1A",X"F3",X"01",X"DC",X"3E",X"A8",X"02",X"B5",X"4B",X"3E",X"62",X"5C",X"DE",
		X"3E",X"62",X"F4",X"00",X"ED",X"0B",X"DC",X"3E",X"3E",X"B6",X"57",X"DE",X"3E",X"62",X"7A",X"63",
		X"33",X"DC",X"3E",X"A8",X"B5",X"76",X"5F",X"60",X"19",X"05",X"ED",X"06",X"76",X"91",X"60",X"7A",
		X"68",X"33",X"76",X"91",X"60",X"71",X"04",X"C0",X"71",X"0E",X"00",X"7A",X"ED",X"33",X"FF",X"D9",
		X"76",X"6E",X"60",X"4B",X"65",X"60",X"F4",X"00",X"ED",X"05",X"D9",X"D1",X"00",X"1A",X"03",X"D9",
		X"D1",X"01",X"B5",X"76",X"E7",X"D0",X"A4",X"25",X"34",X"A4",X"00",X"22",X"B5",X"C0",X"71",X"10",
		X"C0",X"71",X"02",X"C0",X"71",X"03",X"C0",X"71",X"00",X"C0",X"71",X"08",X"C0",X"71",X"01",X"C0",
		X"71",X"0C",X"C0",X"71",X"09",X"C0",X"71",X"0F",X"C0",X"71",X"0A",X"B5",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"D4",X"00",X"25",X"33",X"15",X"00",X"04",X"B3",X"0A",X"CB",X"B3",
		X"0A",X"F8",X"66",X"40",X"08",X"3E",X"C0",X"C0",X"89",X"F7",X"26",X"15",X"2C",X"00",X"40",X"D3",
		X"DC",X"89",X"EB",X"B5",X"04",X"00",X"B5",X"3F",X"7D",X"5E",X"F4",X"64",X"7D",X"5A",X"F4",X"07",
		X"2C",X"24",X"F4",X"09",X"7D",X"20",X"F4",X"31",X"7D",X"1C",X"F4",X"3A",X"7D",X"18",X"F4",X"3C",
		X"7D",X"14",X"F4",X"43",X"7D",X"10",X"F4",X"5A",X"7D",X"0C",X"F4",X"6B",X"7D",X"08",X"F4",X"6D",
		X"7D",X"04",X"F4",X"6E",X"ED",X"03",X"77",X"1A",X"2E",X"F4",X"18",X"7D",X"28",X"F4",X"1C",X"7D",
		X"24",X"F4",X"2C",X"7D",X"20",X"F4",X"3A",X"7D",X"1C",X"F4",X"3B",X"7D",X"18",X"F4",X"3E",X"7D",
		X"14",X"F4",X"56",X"7D",X"10",X"F4",X"6A",X"7D",X"0C",X"F4",X"6C",X"7D",X"08",X"F4",X"6F",X"7D",
		X"04",X"F4",X"70",X"ED",X"02",X"77",X"77",X"77",X"B5",X"A4",X"26",X"1F",X"F4",X"01",X"ED",X"04",
		X"25",X"02",X"1A",X"1A",X"F4",X"05",X"EA",X"04",X"25",X"03",X"1A",X"12",X"F4",X"0A",X"EA",X"04",
		X"25",X"04",X"1A",X"0A",X"F4",X"11",X"EA",X"04",X"25",X"05",X"1A",X"02",X"25",X"06",X"B5",X"FF",
		X"66",X"26",X"CB",X"76",X"AB",X"62",X"4B",X"65",X"60",X"5F",X"ED",X"09",X"19",X"3C",X"ED",X"29",
		X"15",X"66",X"60",X"1A",X"07",X"19",X"FA",X"ED",X"20",X"15",X"67",X"60",X"4B",X"02",X"90",X"6D",
		X"04",X"25",X"02",X"ED",X"02",X"25",X"03",X"D9",X"21",X"00",X"ED",X"0D",X"19",X"5A",X"7B",X"5C",
		X"18",X"76",X"01",X"60",X"19",X"54",X"A4",X"77",X"1D",X"DC",X"D3",X"3E",X"A4",X"06",X"1E",X"B5",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"A4",X"26",X"1F",X"76",X"AA",X"60",X"7A",X"7E",X"22",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"F4",X"06",X"EA",X"04",X"71",X"04",X"1A",X"02",X"71",X"02",X"22",X"C0",X"F8",X"B5",X"76",
		X"5F",X"60",X"19",X"05",X"9B",X"29",X"36",X"45",X"D8",X"61",X"4B",X"27",X"60",X"6D",X"0F",X"F4",
		X"08",X"ED",X"13",X"4B",X"28",X"60",X"6D",X"0F",X"F4",X"06",X"ED",X"0A",X"C0",X"22",X"F4",X"FF",
		X"ED",X"01",X"0C",X"37",X"D8",X"61",X"22",X"1A",X"17",X"4B",X"65",X"60",X"F4",X"00",X"7D",X"0C",
		X"4B",X"02",X"90",X"19",X"EB",X"7D",X"05",X"4B",X"01",X"90",X"1A",X"03",X"4B",X"00",X"90",X"8B",
		X"6D",X"0F",X"31",X"F4",X"01",X"7D",X"0B",X"F4",X"02",X"7D",X"07",X"F4",X"04",X"7D",X"03",X"F4",
		X"08",X"F9",X"48",X"4B",X"5F",X"60",X"19",X"B8",X"9B",X"C1",X"36",X"4B",X"27",X"60",X"6D",X"0F",
		X"F4",X"08",X"9B",X"43",X"49",X"4B",X"28",X"60",X"6D",X"0F",X"F4",X"06",X"F3",X"4B",X"49",X"26",
		X"EE",X"DE",X"E0",X"61",X"7A",X"CE",X"36",X"19",X"02",X"DD",X"F3",X"1E",X"38",X"76",X"27",X"60",
		X"6D",X"0A",X"7D",X"1E",X"22",X"6D",X"0F",X"F4",X"08",X"2C",X"03",X"9E",X"1A",X"01",X"D1",X"C0",
		X"19",X"E8",X"ED",X"07",X"9E",X"25",X"02",X"DE",X"98",X"61",X"B5",X"D1",X"25",X"08",X"DE",X"98",
		X"61",X"B5",X"C0",X"22",X"6D",X"0F",X"F4",X"07",X"2C",X"03",X"9E",X"1A",X"01",X"D1",X"0C",X"19",
		X"29",X"7D",X"07",X"D1",X"25",X"04",X"DE",X"98",X"61",X"B5",X"9E",X"25",X"01",X"DE",X"98",X"61",
		X"B5",X"26",X"EE",X"DE",X"E0",X"61",X"4B",X"98",X"61",X"6D",X"0A",X"F3",X"6E",X"37",X"4B",X"27",
		X"60",X"72",X"4B",X"28",X"60",X"A4",X"DA",X"36",X"1A",X"1B",X"6E",X"36",X"19",X"02",X"19",X"02",
		X"19",X"02",X"19",X"02",X"19",X"99",X"76",X"E4",X"0D",X"CE",X"00",X"57",X"40",X"69",X"C0",X"0D",
		X"25",X"08",X"D4",X"10",X"B5",X"19",X"4B",X"19",X"9D",X"2C",X"03",X"C8",X"1A",X"F7",X"A4",X"03",
		X"37",X"1A",X"03",X"33",X"02",X"B5",X"7D",X"06",X"2C",X"08",X"19",X"30",X"1A",X"ED",X"E9",X"EB",
		X"1A",X"0D",X"E9",X"19",X"C0",X"19",X"18",X"82",X"19",X"C0",X"19",X"18",X"EA",X"F9",X"EB",X"4B",
		X"27",X"60",X"32",X"D9",X"76",X"96",X"61",X"E0",X"6E",X"06",X"48",X"32",X"DD",X"EA",X"33",X"32",
		X"1D",X"6E",X"02",X"48",X"32",X"DD",X"EA",X"25",X"32",X"92",X"5A",X"06",X"57",X"32",X"4C",X"2C",
		X"17",X"32",X"6A",X"5A",X"02",X"57",X"32",X"4C",X"1C",X"0A",X"38",X"D9",X"1F",X"00",X"66",X"76",
		X"E0",X"61",X"19",X"54",X"3E",X"7A",X"0A",X"38",X"D9",X"1F",X"00",X"1A",X"08",X"D9",X"C1",X"00",
		X"1A",X"EC",X"D9",X"C1",X"00",X"4B",X"28",X"60",X"D9",X"F8",X"01",X"7A",X"06",X"38",X"4B",X"28",
		X"60",X"72",X"4B",X"27",X"60",X"A4",X"7A",X"37",X"1A",X"1B",X"6E",X"08",X"19",X"02",X"19",X"02",
		X"19",X"02",X"19",X"02",X"19",X"99",X"76",X"FA",X"0D",X"CE",X"00",X"57",X"40",X"69",X"C0",X"0D",
		X"25",X"36",X"D4",X"10",X"B5",X"19",X"4B",X"19",X"9D",X"2C",X"03",X"C8",X"1A",X"F7",X"A4",X"03",
		X"37",X"7D",X"06",X"2C",X"08",X"19",X"30",X"1A",X"F2",X"E9",X"EB",X"1A",X"0D",X"E9",X"19",X"C0",
		X"19",X"18",X"82",X"19",X"C0",X"19",X"18",X"EA",X"F9",X"EB",X"4B",X"28",X"60",X"32",X"D9",X"76",
		X"96",X"61",X"E0",X"6E",X"05",X"48",X"32",X"DD",X"EA",X"33",X"32",X"1D",X"6E",X"03",X"48",X"32",
		X"DD",X"EA",X"25",X"32",X"92",X"5A",X"05",X"57",X"32",X"4C",X"2C",X"17",X"32",X"6A",X"5A",X"03",
		X"57",X"32",X"4C",X"1C",X"0A",X"38",X"D9",X"1F",X"01",X"66",X"76",X"E0",X"61",X"19",X"5A",X"3E",
		X"7A",X"0A",X"38",X"D9",X"1F",X"01",X"1A",X"08",X"D9",X"C1",X"01",X"1A",X"EC",X"D9",X"C1",X"01",
		X"4B",X"27",X"60",X"D9",X"F8",X"00",X"D3",X"7A",X"8C",X"38",X"D3",X"76",X"5F",X"60",X"19",X"21",
		X"4B",X"26",X"60",X"19",X"02",X"19",X"02",X"19",X"02",X"19",X"02",X"DD",X"7D",X"0F",X"1D",X"19",
		X"99",X"19",X"99",X"19",X"99",X"19",X"99",X"FE",X"02",X"DE",X"26",X"60",X"B5",X"25",X"05",X"A0",
		X"7D",X"0A",X"4B",X"98",X"61",X"6D",X"05",X"9B",X"69",X"38",X"1A",X"08",X"4B",X"98",X"61",X"6D",
		X"0A",X"9B",X"69",X"38",X"D9",X"76",X"27",X"60",X"1D",X"F4",X"02",X"2C",X"0B",X"7D",X"0E",X"F4",
		X"04",X"7D",X"0F",X"D9",X"D1",X"01",X"1A",X"0D",X"D9",X"9E",X"00",X"1A",X"08",X"D9",X"9E",X"01",
		X"1A",X"03",X"D9",X"D1",X"00",X"DE",X"98",X"61",X"B5",X"4B",X"E0",X"61",X"F4",X"00",X"31",X"19",
		X"72",X"7D",X"0D",X"76",X"28",X"60",X"4B",X"97",X"61",X"21",X"2C",X"02",X"D1",X"B5",X"9E",X"B5",
		X"76",X"27",X"60",X"4B",X"96",X"61",X"21",X"2C",X"F5",X"7A",X"7C",X"38",X"76",X"5F",X"60",X"19",
		X"F4",X"4B",X"26",X"60",X"19",X"02",X"19",X"02",X"19",X"02",X"19",X"02",X"DD",X"F3",X"1E",X"38",
		X"E2",X"76",X"26",X"60",X"D9",X"76",X"96",X"61",X"4B",X"28",X"60",X"D9",X"21",X"01",X"ED",X"36",
		X"4B",X"27",X"60",X"D9",X"21",X"00",X"ED",X"07",X"A4",X"0D",X"39",X"1C",X"44",X"38",X"B5",X"4B",
		X"27",X"60",X"D9",X"21",X"00",X"2C",X"10",X"25",X"05",X"A0",X"F3",X"44",X"38",X"A4",X"0D",X"39",
		X"84",X"E2",X"9E",X"01",X"7A",X"44",X"38",X"25",X"05",X"A0",X"ED",X"F8",X"A4",X"0D",X"39",X"84",
		X"E2",X"D1",X"01",X"7A",X"D4",X"38",X"E2",X"22",X"02",X"D9",X"21",X"01",X"2C",X"0F",X"25",X"0A",
		X"A0",X"ED",X"E1",X"A4",X"0D",X"39",X"84",X"E2",X"9E",X"02",X"7A",X"D4",X"38",X"25",X"0A",X"A0",
		X"ED",X"D2",X"A4",X"0D",X"39",X"84",X"E2",X"D1",X"02",X"7A",X"D4",X"38",X"B5",X"D9",X"76",X"96",
		X"61",X"D9",X"22",X"00",X"19",X"02",X"19",X"02",X"19",X"02",X"19",X"02",X"19",X"99",X"57",X"19",
		X"99",X"6B",X"B3",X"00",X"04",X"76",X"A2",X"0D",X"D6",X"D9",X"22",X"01",X"19",X"02",X"19",X"02",
		X"19",X"02",X"19",X"02",X"6E",X"03",X"57",X"19",X"02",X"04",X"D6",X"22",X"19",X"8D",X"7D",X"0B",
		X"19",X"02",X"19",X"02",X"19",X"02",X"19",X"02",X"7A",X"4D",X"39",X"6D",X"0F",X"57",X"A0",X"F3",
		X"54",X"39",X"A8",X"B5",X"0A",X"B5",X"45",X"99",X"61",X"C0",X"37",X"99",X"61",X"92",X"6D",X"08",
		X"F4",X"08",X"25",X"01",X"7D",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"02",X"B3",X"06",X"D9",X"76",X"A8",X"61",X"15",X"00",
		X"04",X"D9",X"24",X"00",X"D9",X"C0",X"D9",X"05",X"00",X"D9",X"C0",X"04",X"EE",X"16",X"C2",X"7D",
		X"0D",X"40",X"F8",X"C0",X"F8",X"26",X"15",X"E0",X"FF",X"40",X"D3",X"F8",X"0C",X"F8",X"89",X"E1",
		X"B5",X"76",X"AA",X"60",X"9E",X"F3",X"48",X"3A",X"76",X"63",X"60",X"9E",X"ED",X"07",X"71",X"03",
		X"76",X"00",X"60",X"19",X"6D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"61",X"60",X"D1",X"22",X"F4",X"17",X"ED",X"0F",
		X"71",X"00",X"76",X"60",X"60",X"D1",X"22",X"F4",X"04",X"ED",X"16",X"71",X"00",X"1A",X"12",X"F4",
		X"0C",X"ED",X"0E",X"4B",X"60",X"60",X"F4",X"00",X"ED",X"07",X"4B",X"62",X"60",X"8B",X"DE",X"62",
		X"60",X"4B",X"AB",X"60",X"DE",X"AA",X"60",X"4B",X"60",X"60",X"F4",X"00",X"ED",X"3A",X"4B",X"61",
		X"60",X"F4",X"01",X"7D",X"1B",X"F4",X"0C",X"ED",X"2F",X"B3",X"04",X"15",X"05",X"00",X"A4",X"A8",
		X"30",X"19",X"3C",X"ED",X"05",X"40",X"89",X"F9",X"1A",X"1E",X"19",X"03",X"19",X"54",X"1A",X"18",
		X"B3",X"04",X"15",X"05",X"00",X"76",X"2B",X"60",X"19",X"3C",X"ED",X"05",X"40",X"89",X"F9",X"1A",
		X"07",X"66",X"76",X"00",X"60",X"19",X"55",X"3E",X"76",X"CA",X"61",X"9E",X"76",X"B6",X"61",X"9E",
		X"C0",X"ED",X"22",X"0C",X"71",X"3C",X"C0",X"66",X"C0",X"D1",X"B3",X"04",X"76",X"CE",X"61",X"EE",
		X"21",X"7D",X"01",X"9E",X"C0",X"89",X"F9",X"76",X"E1",X"61",X"21",X"7D",X"01",X"9E",X"3E",X"22",
		X"F4",X"F0",X"EA",X"01",X"D1",X"C0",X"C0",X"9E",X"B5",X"66",X"26",X"97",X"1D",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"76",X"7A",X"0D",
		X"01",X"57",X"CE",X"00",X"40",X"22",X"D3",X"3E",X"B5",X"4B",X"C9",X"61",X"6D",X"FF",X"7D",X"03",
		X"7A",X"F9",X"3A",X"4B",X"26",X"60",X"19",X"02",X"19",X"02",X"19",X"02",X"19",X"02",X"76",X"98",
		X"61",X"21",X"F9",X"F4",X"02",X"E7",X"98",X"3B",X"9B",X"61",X"3B",X"F4",X"04",X"9B",X"2E",X"3B",
		X"4B",X"27",X"60",X"6E",X"04",X"48",X"4B",X"28",X"60",X"00",X"57",X"A4",X"0A",X"3C",X"3C",X"38",
		X"A4",X"0A",X"3C",X"22",X"33",X"7D",X"21",X"65",X"F4",X"36",X"ED",X"05",X"C0",X"EE",X"7A",X"CA",
		X"3B",X"7C",X"1D",X"5A",X"08",X"48",X"A4",X"0A",X"3C",X"25",X"35",X"21",X"F9",X"26",X"15",X"20",
		X"00",X"40",X"D3",X"25",X"01",X"7A",X"CA",X"3B",X"B5",X"45",X"CB",X"61",X"4B",X"C9",X"61",X"32",
		X"EE",X"DE",X"C9",X"61",X"32",X"F4",X"02",X"7D",X"0A",X"2C",X"0C",X"F4",X"03",X"7D",X"0C",X"25",
		X"06",X"1A",X"0A",X"25",X"07",X"1A",X"06",X"25",X"05",X"1A",X"02",X"25",X"04",X"A4",X"EA",X"3B",
		X"A4",X"EB",X"22",X"A4",X"7B",X"46",X"76",X"5F",X"60",X"19",X"12",X"7A",X"A3",X"3A",X"4B",X"27",
		X"60",X"5A",X"05",X"48",X"4B",X"28",X"60",X"5A",X"05",X"57",X"A4",X"0A",X"3C",X"22",X"78",X"A4",
		X"0A",X"3C",X"21",X"7D",X"1B",X"25",X"3E",X"21",X"ED",X"05",X"25",X"03",X"7A",X"CA",X"3B",X"6A",
		X"6E",X"08",X"57",X"A4",X"0A",X"3C",X"25",X"3D",X"21",X"F9",X"0C",X"25",X"02",X"7A",X"CA",X"3B",
		X"B5",X"4B",X"27",X"60",X"5A",X"04",X"48",X"4B",X"28",X"60",X"6E",X"04",X"57",X"A4",X"0A",X"3C",
		X"22",X"38",X"A4",X"0A",X"3C",X"21",X"7D",X"1F",X"25",X"35",X"21",X"ED",X"0A",X"26",X"15",X"20",
		X"00",X"40",X"D3",X"EE",X"7A",X"CA",X"3B",X"1D",X"6E",X"08",X"48",X"A4",X"0A",X"3C",X"25",X"36",
		X"21",X"F9",X"25",X"01",X"7A",X"CA",X"3B",X"B5",X"7A",X"80",X"00",X"5C",X"48",X"4B",X"28",X"60",
		X"6E",X"03",X"57",X"A4",X"0A",X"3C",X"22",X"2A",X"A4",X"0A",X"3C",X"21",X"7D",X"1B",X"25",X"3D",
		X"21",X"ED",X"06",X"0C",X"25",X"03",X"7A",X"CA",X"3B",X"6A",X"5A",X"08",X"57",X"A4",X"0A",X"3C",
		X"25",X"3E",X"21",X"F9",X"25",X"02",X"7A",X"CA",X"3B",X"B5",X"32",X"4B",X"C9",X"61",X"F4",X"00",
		X"F3",X"F9",X"3A",X"32",X"72",X"5C",X"DE",X"C9",X"61",X"65",X"37",X"CB",X"61",X"32",X"25",X"01",
		X"DE",X"CA",X"61",X"32",X"A4",X"EA",X"3B",X"7A",X"FE",X"3B",X"7A",X"8A",X"56",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"A4",X"EB",
		X"22",X"A4",X"7B",X"46",X"76",X"5F",X"60",X"19",X"12",X"B5",X"97",X"CB",X"1D",X"6D",X"F8",X"B3",
		X"00",X"04",X"19",X"76",X"19",X"89",X"19",X"76",X"19",X"89",X"76",X"A0",X"D0",X"D6",X"6A",X"19",
		X"02",X"19",X"02",X"19",X"02",X"B3",X"00",X"04",X"D6",X"DC",X"01",X"B5",X"66",X"76",X"5F",X"60",
		X"19",X"05",X"F3",X"AE",X"3C",X"26",X"4B",X"65",X"60",X"F4",X"00",X"ED",X"05",X"4B",X"9F",X"60",
		X"1A",X"03",X"4B",X"A2",X"60",X"32",X"76",X"10",X"0E",X"EE",X"4C",X"ED",X"15",X"32",X"B3",X"00",
		X"04",X"D6",X"22",X"19",X"99",X"19",X"99",X"19",X"99",X"19",X"99",X"B3",X"00",X"D4",X"00",X"48",
		X"1A",X"10",X"38",X"19",X"C0",X"19",X"C0",X"CE",X"00",X"40",X"32",X"57",X"40",X"B3",X"00",X"FA",
		X"CE",X"00",X"4B",X"65",X"60",X"F4",X"00",X"ED",X"06",X"D9",X"76",X"68",X"60",X"1A",X"04",X"D9",
		X"76",X"6B",X"60",X"D9",X"22",X"02",X"EC",X"99",X"D9",X"F8",X"02",X"D9",X"22",X"01",X"C3",X"99",
		X"D9",X"F8",X"01",X"D9",X"22",X"00",X"56",X"99",X"D9",X"F8",X"00",X"4B",X"65",X"60",X"F4",X"00",
		X"ED",X"05",X"76",X"C4",X"D2",X"1A",X"03",X"76",X"C3",X"D2",X"A4",X"D0",X"34",X"D3",X"3E",X"B5",
		X"66",X"26",X"CB",X"76",X"44",X"60",X"15",X"FB",X"FF",X"B3",X"06",X"EE",X"19",X"FA",X"7D",X"04",
		X"A8",X"7A",X"C5",X"3C",X"0A",X"BA",X"40",X"89",X"F3",X"DC",X"D3",X"3E",X"B5",X"CB",X"26",X"66",
		X"B3",X"09",X"15",X"05",X"00",X"76",X"21",X"60",X"19",X"03",X"19",X"4A",X"40",X"89",X"F9",X"D9",
		X"66",X"E2",X"66",X"97",X"A4",X"C7",X"1F",X"A4",X"8F",X"17",X"01",X"E2",X"3E",X"D9",X"3E",X"3E",
		X"D3",X"DC",X"B5",X"D9",X"76",X"43",X"0D",X"B3",X"14",X"F2",X"00",X"D9",X"24",X"00",X"D9",X"05",
		X"01",X"22",X"F4",X"36",X"ED",X"03",X"0A",X"1A",X"01",X"A8",X"19",X"C7",X"19",X"18",X"19",X"15",
		X"D9",X"0C",X"D9",X"0C",X"89",X"E5",X"4B",X"65",X"60",X"F4",X"00",X"ED",X"05",X"76",X"A3",X"60",
		X"1A",X"03",X"76",X"A6",X"60",X"07",X"C0",X"91",X"C0",X"08",X"B5",X"66",X"D4",X"02",X"B3",X"03",
		X"15",X"02",X"0C",X"7B",X"C7",X"3A",X"F3",X"3E",X"3D",X"7B",X"16",X"9B",X"64",X"3D",X"C7",X"89",
		X"F2",X"9A",X"B3",X"03",X"7B",X"C7",X"3A",X"F3",X"4F",X"3D",X"7B",X"16",X"9B",X"64",X"3D",X"C7",
		X"89",X"F2",X"D4",X"03",X"00",X"7A",X"64",X"3D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B3",X"00",X"D9",X"76",X"58",X"0E",X"19",X"76",X"19",X"76",X"D9",X"D6",
		X"D9",X"22",X"00",X"F8",X"66",X"15",X"00",X"04",X"40",X"71",X"02",X"3E",X"C0",X"D9",X"22",X"01",
		X"F8",X"66",X"40",X"71",X"00",X"3E",X"26",X"15",X"E0",X"FF",X"40",X"D3",X"D9",X"22",X"02",X"F8",
		X"66",X"40",X"71",X"00",X"3E",X"0C",X"D9",X"22",X"03",X"F8",X"40",X"71",X"00",X"3E",X"B5",X"66",
		X"45",X"99",X"61",X"E0",X"F4",X"00",X"ED",X"09",X"92",X"F4",X"1F",X"2C",X"08",X"F4",X"B4",X"2C",
		X"08",X"F2",X"01",X"1A",X"06",X"F2",X"03",X"1A",X"02",X"F2",X"02",X"3E",X"B5",X"26",X"25",X"DA",
		X"32",X"4B",X"65",X"60",X"F4",X"00",X"ED",X"05",X"4B",X"9F",X"60",X"1A",X"03",X"4B",X"A2",X"60",
		X"F4",X"00",X"7D",X"0D",X"F4",X"03",X"7D",X"06",X"72",X"32",X"23",X"17",X"1A",X"02",X"25",X"DD",
		X"F8",X"D9",X"76",X"26",X"60",X"D9",X"19",X"00",X"86",X"D9",X"19",X"00",X"8E",X"D9",X"76",X"49",
		X"60",X"D9",X"71",X"00",X"82",X"7A",X"F0",X"2F",X"25",X"09",X"C8",X"D9",X"F8",X"02",X"D9",X"A3",
		X"01",X"D9",X"71",X"04",X"03",X"6A",X"F4",X"02",X"2C",X"0E",X"7D",X"06",X"D9",X"71",X"03",X"E0",
		X"1A",X"0A",X"D9",X"71",X"03",X"DC",X"1A",X"04",X"D9",X"71",X"03",X"D8",X"66",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A4",X"4A",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"EE",X"DE",X"49",X"60",X"76",X"26",X"60",X"19",X"54",X"3E",X"71",X"FF",X"D3",X"B5",X"66",
		X"26",X"15",X"A0",X"D0",X"0A",X"B6",X"29",X"47",X"25",X"E0",X"E5",X"EB",X"B3",X"02",X"19",X"5C",
		X"19",X"38",X"89",X"FA",X"43",X"19",X"76",X"19",X"76",X"19",X"76",X"D3",X"3E",X"B5",X"66",X"CE",
		X"00",X"F4",X"5E",X"7D",X"2F",X"78",X"F4",X"5B",X"7D",X"2A",X"78",X"F4",X"59",X"7D",X"25",X"78",
		X"F4",X"5A",X"7D",X"20",X"78",X"F4",X"5C",X"ED",X"0A",X"C0",X"22",X"F4",X"66",X"2C",X"15",X"78",
		X"78",X"1A",X"11",X"78",X"F4",X"5D",X"7D",X"0C",X"78",X"78",X"F4",X"5F",X"7D",X"06",X"78",X"F4",
		X"60",X"7D",X"01",X"78",X"3E",X"B5",X"F4",X"03",X"7D",X"05",X"F4",X"02",X"7D",X"12",X"B5",X"4B",
		X"65",X"60",X"F4",X"00",X"ED",X"05",X"76",X"9D",X"60",X"1A",X"16",X"76",X"A0",X"60",X"1A",X"11",
		X"4B",X"65",X"60",X"F4",X"00",X"ED",X"05",X"76",X"9E",X"60",X"1A",X"3E",X"76",X"A1",X"60",X"1A",
		X"39",X"1D",X"F4",X"00",X"ED",X"04",X"19",X"AA",X"1A",X"2E",X"F4",X"01",X"ED",X"04",X"19",X"AC",
		X"1A",X"26",X"F4",X"02",X"ED",X"04",X"19",X"03",X"1A",X"1E",X"F4",X"03",X"ED",X"04",X"19",X"4A",
		X"1A",X"16",X"F4",X"04",X"ED",X"04",X"19",X"12",X"1A",X"0E",X"F4",X"05",X"ED",X"04",X"19",X"CD",
		X"1A",X"06",X"F4",X"06",X"ED",X"02",X"19",X"11",X"1A",X"2F",X"1D",X"F4",X"00",X"ED",X"04",X"19",
		X"CD",X"1A",X"1E",X"F4",X"01",X"ED",X"04",X"19",X"03",X"1A",X"16",X"F4",X"07",X"ED",X"04",X"19",
		X"4A",X"1A",X"0E",X"F4",X"08",X"ED",X"04",X"19",X"AC",X"1A",X"06",X"F4",X"09",X"ED",X"02",X"19",
		X"12",X"0C",X"66",X"A4",X"1C",X"31",X"3E",X"1A",X"05",X"66",X"A4",X"F4",X"30",X"3E",X"B5",X"A4",
		X"C7",X"1F",X"A4",X"8F",X"17",X"4B",X"03",X"60",X"F4",X"00",X"ED",X"F3",X"B5",X"E2",X"76",X"9C",
		X"61",X"D9",X"76",X"91",X"60",X"A4",X"35",X"40",X"D9",X"76",X"92",X"60",X"A4",X"35",X"40",X"D9",
		X"76",X"93",X"60",X"A4",X"35",X"40",X"D9",X"76",X"94",X"60",X"A4",X"35",X"40",X"B5",X"F5",X"D1",
		X"32",X"72",X"25",X"06",X"49",X"7D",X"13",X"72",X"32",X"19",X"99",X"CE",X"00",X"57",X"76",X"A8",
		X"61",X"40",X"71",X"00",X"C0",X"71",X"00",X"C0",X"89",X"F8",X"B5",X"D9",X"66",X"97",X"26",X"65",
		X"F4",X"0A",X"2C",X"12",X"7D",X"0A",X"F4",X"0B",X"ED",X"2D",X"D9",X"76",X"A8",X"61",X"1A",X"0A",
		X"D9",X"76",X"A2",X"61",X"1A",X"04",X"D9",X"76",X"9C",X"61",X"D9",X"22",X"01",X"F4",X"00",X"7D",
		X"10",X"D9",X"C0",X"D9",X"C0",X"D9",X"66",X"15",X"B4",X"61",X"6A",X"D3",X"4C",X"7D",X"08",X"1A",
		X"E9",X"D9",X"1F",X"00",X"D9",X"C1",X"01",X"D3",X"01",X"D9",X"3E",X"B5",X"97",X"CB",X"66",X"EE",
		X"B3",X"18",X"76",X"9C",X"61",X"F8",X"C0",X"89",X"FC",X"3E",X"DC",X"01",X"B5",X"76",X"02",X"90",
		X"19",X"24",X"7D",X"10",X"76",X"00",X"A0",X"4B",X"65",X"60",X"F4",X"00",X"ED",X"04",X"19",X"03",
		X"1A",X"02",X"19",X"5A",X"B5",X"97",X"CB",X"26",X"B3",X"0C",X"15",X"9C",X"61",X"7B",X"3A",X"ED",
		X"06",X"C7",X"7B",X"9D",X"16",X"7D",X"06",X"C7",X"C7",X"89",X"F2",X"1A",X"04",X"EE",X"18",X"C7");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
